entity wifi_tele_logic is

end entity;


architecture arch of wifi_tele_logic is

begin

end arch;