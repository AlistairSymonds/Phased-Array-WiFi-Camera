-- WiPhase_top_level.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity WiPhase_top_level is
	port (
		mac_mdio_connection_mdc           : out std_logic;                                        --       mac_mdio_connection.mdc
		mac_mdio_connection_mdio_in       : in  std_logic                     := '0';             --                          .mdio_in
		mac_mdio_connection_mdio_out      : out std_logic;                                        --                          .mdio_out
		mac_mdio_connection_mdio_oen      : out std_logic;                                        --                          .mdio_oen
		mac_misc_connection_ff_tx_crc_fwd : in  std_logic                     := '0';             --       mac_misc_connection.ff_tx_crc_fwd
		mac_misc_connection_ff_tx_septy   : out std_logic;                                        --                          .ff_tx_septy
		mac_misc_connection_tx_ff_uflow   : out std_logic;                                        --                          .tx_ff_uflow
		mac_misc_connection_ff_tx_a_full  : out std_logic;                                        --                          .ff_tx_a_full
		mac_misc_connection_ff_tx_a_empty : out std_logic;                                        --                          .ff_tx_a_empty
		mac_misc_connection_rx_err_stat   : out std_logic_vector(17 downto 0);                    --                          .rx_err_stat
		mac_misc_connection_rx_frm_type   : out std_logic_vector(3 downto 0);                     --                          .rx_frm_type
		mac_misc_connection_ff_rx_dsav    : out std_logic;                                        --                          .ff_rx_dsav
		mac_misc_connection_ff_rx_a_full  : out std_logic;                                        --                          .ff_rx_a_full
		mac_misc_connection_ff_rx_a_empty : out std_logic;                                        --                          .ff_rx_a_empty
		mac_status_set_10                 : in  std_logic                     := '0';             --                mac_status.set_10
		mac_status_set_1000               : in  std_logic                     := '0';             --                          .set_1000
		mac_status_eth_mode               : out std_logic;                                        --                          .eth_mode
		mac_status_ena_10                 : out std_logic;                                        --                          .ena_10
		mclk_i_clk                        : in  std_logic                     := '0';             --                    mclk_i.clk
		mclk_reset_reset_n                : in  std_logic                     := '0';             --                mclk_reset.reset_n
		pll_inclk_clk                     : in  std_logic                     := '0';             --                 pll_inclk.clk
		pll_out_clk                       : out std_logic;                                        --                   pll_out.clk
		rgmii_connection_rgmii_in         : in  std_logic_vector(3 downto 0)  := (others => '0'); --          rgmii_connection.rgmii_in
		rgmii_connection_rgmii_out        : out std_logic_vector(3 downto 0);                     --                          .rgmii_out
		rgmii_connection_rx_control       : in  std_logic                     := '0';             --                          .rx_control
		rgmii_connection_tx_control       : out std_logic;                                        --                          .tx_control
		rgmii_rx_clk_clk                  : in  std_logic                     := '0';             --              rgmii_rx_clk.clk
		rgmii_tx_clk_clk                  : in  std_logic                     := '0';             --              rgmii_tx_clk.clk
		sample_pll_areset_conduit_export  : in  std_logic                     := '0';             -- sample_pll_areset_conduit.export
		sample_pll_locked_conduit_export  : out std_logic;                                        -- sample_pll_locked_conduit.export
		spi_signals_o_MISO                : in  std_logic                     := '0';             --             spi_signals_o.MISO
		spi_signals_o_MOSI                : out std_logic;                                        --                          .MOSI
		spi_signals_o_SCLK                : out std_logic;                                        --                          .SCLK
		spi_signals_o_SS_n                : out std_logic_vector(2 downto 0)                      --                          .SS_n
	);
end entity WiPhase_top_level;

architecture rtl of WiPhase_top_level is
	component Debug_ST_Sink is
		port (
			ST_sink_connection_data          : in std_logic_vector(7 downto 0) := (others => 'X'); -- data
			ST_sink_connection_endofpacket   : in std_logic                    := 'X';             -- endofpacket
			ST_sink_connection_startofpacket : in std_logic                    := 'X';             -- startofpacket
			clk                              : in std_logic                    := 'X'              -- clk
		);
	end component Debug_ST_Sink;

	component WiPhase_top_level_cpu_v2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(16 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(16 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component WiPhase_top_level_cpu_v2;

	component WiPhase_top_level_eth is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			reg_addr      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			reg_data_out  : out std_logic_vector(31 downto 0);                    -- readdata
			reg_rd        : in  std_logic                     := 'X';             -- read
			reg_data_in   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reg_wr        : in  std_logic                     := 'X';             -- write
			reg_busy      : out std_logic;                                        -- waitrequest
			tx_clk        : in  std_logic                     := 'X';             -- clk
			rx_clk        : in  std_logic                     := 'X';             -- clk
			set_10        : in  std_logic                     := 'X';             -- set_10
			set_1000      : in  std_logic                     := 'X';             -- set_1000
			eth_mode      : out std_logic;                                        -- eth_mode
			ena_10        : out std_logic;                                        -- ena_10
			rgmii_in      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- rgmii_in
			rgmii_out     : out std_logic_vector(3 downto 0);                     -- rgmii_out
			rx_control    : in  std_logic                     := 'X';             -- rx_control
			tx_control    : out std_logic;                                        -- tx_control
			ff_rx_clk     : in  std_logic                     := 'X';             -- clk
			ff_tx_clk     : in  std_logic                     := 'X';             -- clk
			ff_rx_data    : out std_logic_vector(31 downto 0);                    -- data
			ff_rx_eop     : out std_logic;                                        -- endofpacket
			rx_err        : out std_logic_vector(5 downto 0);                     -- error
			ff_rx_mod     : out std_logic_vector(1 downto 0);                     -- empty
			ff_rx_rdy     : in  std_logic                     := 'X';             -- ready
			ff_rx_sop     : out std_logic;                                        -- startofpacket
			ff_rx_dval    : out std_logic;                                        -- valid
			ff_tx_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			ff_tx_eop     : in  std_logic                     := 'X';             -- endofpacket
			ff_tx_err     : in  std_logic                     := 'X';             -- error
			ff_tx_mod     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			ff_tx_rdy     : out std_logic;                                        -- ready
			ff_tx_sop     : in  std_logic                     := 'X';             -- startofpacket
			ff_tx_wren    : in  std_logic                     := 'X';             -- valid
			mdc           : out std_logic;                                        -- mdc
			mdio_in       : in  std_logic                     := 'X';             -- mdio_in
			mdio_out      : out std_logic;                                        -- mdio_out
			mdio_oen      : out std_logic;                                        -- mdio_oen
			ff_tx_crc_fwd : in  std_logic                     := 'X';             -- ff_tx_crc_fwd
			ff_tx_septy   : out std_logic;                                        -- ff_tx_septy
			tx_ff_uflow   : out std_logic;                                        -- tx_ff_uflow
			ff_tx_a_full  : out std_logic;                                        -- ff_tx_a_full
			ff_tx_a_empty : out std_logic;                                        -- ff_tx_a_empty
			rx_err_stat   : out std_logic_vector(17 downto 0);                    -- rx_err_stat
			rx_frm_type   : out std_logic_vector(3 downto 0);                     -- rx_frm_type
			ff_rx_dsav    : out std_logic;                                        -- ff_rx_dsav
			ff_rx_a_full  : out std_logic;                                        -- ff_rx_a_full
			ff_rx_a_empty : out std_logic                                         -- ff_rx_a_empty
		);
	end component WiPhase_top_level_eth;

	component WiPhase_top_level_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component WiPhase_top_level_jtag_uart;

	component WiPhase_top_level_ram_onchip is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component WiPhase_top_level_ram_onchip;

	component WiPhase_top_level_sample_pll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			inclk0             : in  std_logic                     := 'X';             -- clk
			c0                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component WiPhase_top_level_sample_pll;

	component WiPhase_top_level_spi is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic_vector(2 downto 0)                      -- export
		);
	end component WiPhase_top_level_spi;

	component WiPhase_top_level_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component WiPhase_top_level_sysid;

	component WiPhase_top_level_test_pattern_st_gen is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset_n             : in  std_logic                     := 'X';             -- reset_n
			csr_address         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_writedata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			csr_read            : in  std_logic                     := 'X';             -- read
			csr_write           : in  std_logic                     := 'X';             -- write
			csr_waitrequest     : out std_logic;                                        -- waitrequest
			command_address     : in  std_logic                     := 'X';             -- address
			command_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			command_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			command_read        : in  std_logic                     := 'X';             -- read
			command_write       : in  std_logic                     := 'X';             -- write
			command_waitrequest : out std_logic;                                        -- waitrequest
			out_valid           : out std_logic;                                        -- valid
			out_data            : out std_logic_vector(7 downto 0);                     -- data
			out_ready           : in  std_logic                     := 'X';             -- ready
			out_startofpacket   : out std_logic;                                        -- startofpacket
			out_endofpacket     : out std_logic                                         -- endofpacket
		);
	end component WiPhase_top_level_test_pattern_st_gen;

	component WiPhase_top_level_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component WiPhase_top_level_timer;

	component WiPhase_top_level_mm_interconnect_0 is
		port (
			C10_Clk50M_clk_clk                       : in  std_logic                     := 'X';             -- clk
			cpu_v2_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_v2_data_master_address               : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			cpu_v2_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			cpu_v2_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_v2_data_master_read                  : in  std_logic                     := 'X';             -- read
			cpu_v2_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_v2_data_master_write                 : in  std_logic                     := 'X';             -- write
			cpu_v2_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_v2_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			cpu_v2_instruction_master_address        : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			cpu_v2_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			cpu_v2_instruction_master_read           : in  std_logic                     := 'X';             -- read
			cpu_v2_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_v2_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			cpu_v2_debug_mem_slave_write             : out std_logic;                                        -- write
			cpu_v2_debug_mem_slave_read              : out std_logic;                                        -- read
			cpu_v2_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_v2_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_v2_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_v2_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			cpu_v2_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			eth_control_port_address                 : out std_logic_vector(7 downto 0);                     -- address
			eth_control_port_write                   : out std_logic;                                        -- write
			eth_control_port_read                    : out std_logic;                                        -- read
			eth_control_port_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			eth_control_port_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			eth_control_port_waitrequest             : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_address      : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write        : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read         : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect   : out std_logic;                                        -- chipselect
			ram_onchip_s1_address                    : out std_logic_vector(12 downto 0);                    -- address
			ram_onchip_s1_write                      : out std_logic;                                        -- write
			ram_onchip_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ram_onchip_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			ram_onchip_s1_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			ram_onchip_s1_chipselect                 : out std_logic;                                        -- chipselect
			ram_onchip_s1_clken                      : out std_logic;                                        -- clken
			sample_pll_pll_slave_address             : out std_logic_vector(1 downto 0);                     -- address
			sample_pll_pll_slave_write               : out std_logic;                                        -- write
			sample_pll_pll_slave_read                : out std_logic;                                        -- read
			sample_pll_pll_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sample_pll_pll_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			spi_spi_control_port_address             : out std_logic_vector(2 downto 0);                     -- address
			spi_spi_control_port_write               : out std_logic;                                        -- write
			spi_spi_control_port_read                : out std_logic;                                        -- read
			spi_spi_control_port_readdata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			spi_spi_control_port_writedata           : out std_logic_vector(15 downto 0);                    -- writedata
			spi_spi_control_port_chipselect          : out std_logic;                                        -- chipselect
			sysid_control_slave_address              : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			test_pattern_st_gen_command_address      : out std_logic_vector(0 downto 0);                     -- address
			test_pattern_st_gen_command_write        : out std_logic;                                        -- write
			test_pattern_st_gen_command_read         : out std_logic;                                        -- read
			test_pattern_st_gen_command_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			test_pattern_st_gen_command_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			test_pattern_st_gen_command_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			test_pattern_st_gen_csr_address          : out std_logic_vector(1 downto 0);                     -- address
			test_pattern_st_gen_csr_write            : out std_logic;                                        -- write
			test_pattern_st_gen_csr_read             : out std_logic;                                        -- read
			test_pattern_st_gen_csr_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			test_pattern_st_gen_csr_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			test_pattern_st_gen_csr_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			timer_s1_address                         : out std_logic_vector(2 downto 0);                     -- address
			timer_s1_write                           : out std_logic;                                        -- write
			timer_s1_readdata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_s1_writedata                       : out std_logic_vector(15 downto 0);                    -- writedata
			timer_s1_chipselect                      : out std_logic                                         -- chipselect
		);
	end component WiPhase_top_level_mm_interconnect_0;

	component WiPhase_top_level_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component WiPhase_top_level_irq_mapper;

	component WiPhase_top_level_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_empty         : out std_logic_vector(1 downto 0);                     -- empty
			out_0_error         : out std_logic_vector(0 downto 0)                      -- error
		);
	end component WiPhase_top_level_avalon_st_adapter;

	component WiPhase_top_level_avalon_st_adapter_001 is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_0_error          : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			out_0_data          : out std_logic_vector(7 downto 0);                     -- data
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component WiPhase_top_level_avalon_st_adapter_001;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal cpu_v2_data_master_readdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_v2_data_master_readdata -> cpu_v2:d_readdata
	signal cpu_v2_data_master_waitrequest                                : std_logic;                     -- mm_interconnect_0:cpu_v2_data_master_waitrequest -> cpu_v2:d_waitrequest
	signal cpu_v2_data_master_debugaccess                                : std_logic;                     -- cpu_v2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_v2_data_master_debugaccess
	signal cpu_v2_data_master_address                                    : std_logic_vector(16 downto 0); -- cpu_v2:d_address -> mm_interconnect_0:cpu_v2_data_master_address
	signal cpu_v2_data_master_byteenable                                 : std_logic_vector(3 downto 0);  -- cpu_v2:d_byteenable -> mm_interconnect_0:cpu_v2_data_master_byteenable
	signal cpu_v2_data_master_read                                       : std_logic;                     -- cpu_v2:d_read -> mm_interconnect_0:cpu_v2_data_master_read
	signal cpu_v2_data_master_write                                      : std_logic;                     -- cpu_v2:d_write -> mm_interconnect_0:cpu_v2_data_master_write
	signal cpu_v2_data_master_writedata                                  : std_logic_vector(31 downto 0); -- cpu_v2:d_writedata -> mm_interconnect_0:cpu_v2_data_master_writedata
	signal cpu_v2_instruction_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_v2_instruction_master_readdata -> cpu_v2:i_readdata
	signal cpu_v2_instruction_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:cpu_v2_instruction_master_waitrequest -> cpu_v2:i_waitrequest
	signal cpu_v2_instruction_master_address                             : std_logic_vector(16 downto 0); -- cpu_v2:i_address -> mm_interconnect_0:cpu_v2_instruction_master_address
	signal cpu_v2_instruction_master_read                                : std_logic;                     -- cpu_v2:i_read -> mm_interconnect_0:cpu_v2_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_test_pattern_st_gen_command_readdata        : std_logic_vector(31 downto 0); -- test_pattern_st_gen:command_readdata -> mm_interconnect_0:test_pattern_st_gen_command_readdata
	signal mm_interconnect_0_test_pattern_st_gen_command_waitrequest     : std_logic;                     -- test_pattern_st_gen:command_waitrequest -> mm_interconnect_0:test_pattern_st_gen_command_waitrequest
	signal mm_interconnect_0_test_pattern_st_gen_command_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:test_pattern_st_gen_command_address -> test_pattern_st_gen:command_address
	signal mm_interconnect_0_test_pattern_st_gen_command_read            : std_logic;                     -- mm_interconnect_0:test_pattern_st_gen_command_read -> test_pattern_st_gen:command_read
	signal mm_interconnect_0_test_pattern_st_gen_command_write           : std_logic;                     -- mm_interconnect_0:test_pattern_st_gen_command_write -> test_pattern_st_gen:command_write
	signal mm_interconnect_0_test_pattern_st_gen_command_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:test_pattern_st_gen_command_writedata -> test_pattern_st_gen:command_writedata
	signal mm_interconnect_0_eth_control_port_readdata                   : std_logic_vector(31 downto 0); -- eth:reg_data_out -> mm_interconnect_0:eth_control_port_readdata
	signal mm_interconnect_0_eth_control_port_waitrequest                : std_logic;                     -- eth:reg_busy -> mm_interconnect_0:eth_control_port_waitrequest
	signal mm_interconnect_0_eth_control_port_address                    : std_logic_vector(7 downto 0);  -- mm_interconnect_0:eth_control_port_address -> eth:reg_addr
	signal mm_interconnect_0_eth_control_port_read                       : std_logic;                     -- mm_interconnect_0:eth_control_port_read -> eth:reg_rd
	signal mm_interconnect_0_eth_control_port_write                      : std_logic;                     -- mm_interconnect_0:eth_control_port_write -> eth:reg_wr
	signal mm_interconnect_0_eth_control_port_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:eth_control_port_writedata -> eth:reg_data_in
	signal mm_interconnect_0_sysid_control_slave_readdata                : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                 : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_test_pattern_st_gen_csr_readdata            : std_logic_vector(31 downto 0); -- test_pattern_st_gen:csr_readdata -> mm_interconnect_0:test_pattern_st_gen_csr_readdata
	signal mm_interconnect_0_test_pattern_st_gen_csr_waitrequest         : std_logic;                     -- test_pattern_st_gen:csr_waitrequest -> mm_interconnect_0:test_pattern_st_gen_csr_waitrequest
	signal mm_interconnect_0_test_pattern_st_gen_csr_address             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:test_pattern_st_gen_csr_address -> test_pattern_st_gen:csr_address
	signal mm_interconnect_0_test_pattern_st_gen_csr_read                : std_logic;                     -- mm_interconnect_0:test_pattern_st_gen_csr_read -> test_pattern_st_gen:csr_read
	signal mm_interconnect_0_test_pattern_st_gen_csr_write               : std_logic;                     -- mm_interconnect_0:test_pattern_st_gen_csr_write -> test_pattern_st_gen:csr_write
	signal mm_interconnect_0_test_pattern_st_gen_csr_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:test_pattern_st_gen_csr_writedata -> test_pattern_st_gen:csr_writedata
	signal mm_interconnect_0_cpu_v2_debug_mem_slave_readdata             : std_logic_vector(31 downto 0); -- cpu_v2:debug_mem_slave_readdata -> mm_interconnect_0:cpu_v2_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_v2_debug_mem_slave_waitrequest          : std_logic;                     -- cpu_v2:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_v2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_v2_debug_mem_slave_debugaccess          : std_logic;                     -- mm_interconnect_0:cpu_v2_debug_mem_slave_debugaccess -> cpu_v2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_v2_debug_mem_slave_address              : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_v2_debug_mem_slave_address -> cpu_v2:debug_mem_slave_address
	signal mm_interconnect_0_cpu_v2_debug_mem_slave_read                 : std_logic;                     -- mm_interconnect_0:cpu_v2_debug_mem_slave_read -> cpu_v2:debug_mem_slave_read
	signal mm_interconnect_0_cpu_v2_debug_mem_slave_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_v2_debug_mem_slave_byteenable -> cpu_v2:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_v2_debug_mem_slave_write                : std_logic;                     -- mm_interconnect_0:cpu_v2_debug_mem_slave_write -> cpu_v2:debug_mem_slave_write
	signal mm_interconnect_0_cpu_v2_debug_mem_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_v2_debug_mem_slave_writedata -> cpu_v2:debug_mem_slave_writedata
	signal mm_interconnect_0_sample_pll_pll_slave_readdata               : std_logic_vector(31 downto 0); -- sample_pll:readdata -> mm_interconnect_0:sample_pll_pll_slave_readdata
	signal mm_interconnect_0_sample_pll_pll_slave_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sample_pll_pll_slave_address -> sample_pll:address
	signal mm_interconnect_0_sample_pll_pll_slave_read                   : std_logic;                     -- mm_interconnect_0:sample_pll_pll_slave_read -> sample_pll:read
	signal mm_interconnect_0_sample_pll_pll_slave_write                  : std_logic;                     -- mm_interconnect_0:sample_pll_pll_slave_write -> sample_pll:write
	signal mm_interconnect_0_sample_pll_pll_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:sample_pll_pll_slave_writedata -> sample_pll:writedata
	signal mm_interconnect_0_ram_onchip_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:ram_onchip_s1_chipselect -> ram_onchip:chipselect
	signal mm_interconnect_0_ram_onchip_s1_readdata                      : std_logic_vector(31 downto 0); -- ram_onchip:readdata -> mm_interconnect_0:ram_onchip_s1_readdata
	signal mm_interconnect_0_ram_onchip_s1_address                       : std_logic_vector(12 downto 0); -- mm_interconnect_0:ram_onchip_s1_address -> ram_onchip:address
	signal mm_interconnect_0_ram_onchip_s1_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ram_onchip_s1_byteenable -> ram_onchip:byteenable
	signal mm_interconnect_0_ram_onchip_s1_write                         : std_logic;                     -- mm_interconnect_0:ram_onchip_s1_write -> ram_onchip:write
	signal mm_interconnect_0_ram_onchip_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:ram_onchip_s1_writedata -> ram_onchip:writedata
	signal mm_interconnect_0_ram_onchip_s1_clken                         : std_logic;                     -- mm_interconnect_0:ram_onchip_s1_clken -> ram_onchip:clken
	signal mm_interconnect_0_timer_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	signal mm_interconnect_0_timer_s1_readdata                           : std_logic_vector(15 downto 0); -- timer:readdata -> mm_interconnect_0:timer_s1_readdata
	signal mm_interconnect_0_timer_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_s1_address -> timer:address
	signal mm_interconnect_0_timer_s1_write                              : std_logic;                     -- mm_interconnect_0:timer_s1_write -> mm_interconnect_0_timer_s1_write:in
	signal mm_interconnect_0_timer_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_s1_writedata -> timer:writedata
	signal mm_interconnect_0_spi_spi_control_port_chipselect             : std_logic;                     -- mm_interconnect_0:spi_spi_control_port_chipselect -> spi:spi_select
	signal mm_interconnect_0_spi_spi_control_port_readdata               : std_logic_vector(15 downto 0); -- spi:data_to_cpu -> mm_interconnect_0:spi_spi_control_port_readdata
	signal mm_interconnect_0_spi_spi_control_port_address                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_spi_control_port_address -> spi:mem_addr
	signal mm_interconnect_0_spi_spi_control_port_read                   : std_logic;                     -- mm_interconnect_0:spi_spi_control_port_read -> mm_interconnect_0_spi_spi_control_port_read:in
	signal mm_interconnect_0_spi_spi_control_port_write                  : std_logic;                     -- mm_interconnect_0:spi_spi_control_port_write -> mm_interconnect_0_spi_spi_control_port_write:in
	signal mm_interconnect_0_spi_spi_control_port_writedata              : std_logic_vector(15 downto 0); -- mm_interconnect_0:spi_spi_control_port_writedata -> spi:data_from_cpu
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- spi:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- timer:irq -> irq_mapper:receiver2_irq
	signal cpu_v2_irq_irq                                                : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu_v2:irq
	signal test_pattern_st_gen_out_valid                                 : std_logic;                     -- test_pattern_st_gen:out_valid -> avalon_st_adapter:in_0_valid
	signal test_pattern_st_gen_out_data                                  : std_logic_vector(7 downto 0);  -- test_pattern_st_gen:out_data -> avalon_st_adapter:in_0_data
	signal test_pattern_st_gen_out_ready                                 : std_logic;                     -- avalon_st_adapter:in_0_ready -> test_pattern_st_gen:out_ready
	signal test_pattern_st_gen_out_startofpacket                         : std_logic;                     -- test_pattern_st_gen:out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	signal test_pattern_st_gen_out_endofpacket                           : std_logic;                     -- test_pattern_st_gen:out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	signal avalon_st_adapter_out_0_valid                                 : std_logic;                     -- avalon_st_adapter:out_0_valid -> eth:ff_tx_wren
	signal avalon_st_adapter_out_0_data                                  : std_logic_vector(31 downto 0); -- avalon_st_adapter:out_0_data -> eth:ff_tx_data
	signal avalon_st_adapter_out_0_ready                                 : std_logic;                     -- eth:ff_tx_rdy -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket                         : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> eth:ff_tx_sop
	signal avalon_st_adapter_out_0_endofpacket                           : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> eth:ff_tx_eop
	signal avalon_st_adapter_out_0_error                                 : std_logic_vector(0 downto 0);  -- avalon_st_adapter:out_0_error -> eth:ff_tx_err
	signal avalon_st_adapter_out_0_empty                                 : std_logic_vector(1 downto 0);  -- avalon_st_adapter:out_0_empty -> eth:ff_tx_mod
	signal eth_receive_valid                                             : std_logic;                     -- eth:ff_rx_dval -> avalon_st_adapter_001:in_0_valid
	signal eth_receive_data                                              : std_logic_vector(31 downto 0); -- eth:ff_rx_data -> avalon_st_adapter_001:in_0_data
	signal eth_receive_ready                                             : std_logic;                     -- avalon_st_adapter_001:in_0_ready -> eth:ff_rx_rdy
	signal eth_receive_startofpacket                                     : std_logic;                     -- eth:ff_rx_sop -> avalon_st_adapter_001:in_0_startofpacket
	signal eth_receive_endofpacket                                       : std_logic;                     -- eth:ff_rx_eop -> avalon_st_adapter_001:in_0_endofpacket
	signal eth_receive_error                                             : std_logic_vector(5 downto 0);  -- eth:rx_err -> avalon_st_adapter_001:in_0_error
	signal eth_receive_empty                                             : std_logic_vector(1 downto 0);  -- eth:ff_rx_mod -> avalon_st_adapter_001:in_0_empty
	signal avalon_st_adapter_001_out_0_data                              : std_logic_vector(7 downto 0);  -- avalon_st_adapter_001:out_0_data -> Debug_ST_Sink_0:ST_sink_connection_data
	signal avalon_st_adapter_001_out_0_startofpacket                     : std_logic;                     -- avalon_st_adapter_001:out_0_startofpacket -> Debug_ST_Sink_0:ST_sink_connection_startofpacket
	signal avalon_st_adapter_001_out_0_endofpacket                       : std_logic;                     -- avalon_st_adapter_001:out_0_endofpacket -> Debug_ST_Sink_0:ST_sink_connection_endofpacket
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, eth:reset, irq_mapper:reset, mm_interconnect_0:cpu_v2_reset_reset_bridge_in_reset_reset, ram_onchip:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, sample_pll:reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [cpu_v2:reset_req, ram_onchip:reset_req, rst_translator:reset_req_in]
	signal mclk_reset_reset_n_ports_inv                                  : std_logic;                     -- mclk_reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_timer_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_timer_s1_write:inv -> timer:write_n
	signal mm_interconnect_0_spi_spi_control_port_read_ports_inv         : std_logic;                     -- mm_interconnect_0_spi_spi_control_port_read:inv -> spi:read_n
	signal mm_interconnect_0_spi_spi_control_port_write_ports_inv        : std_logic;                     -- mm_interconnect_0_spi_spi_control_port_write:inv -> spi:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu_v2:reset_n, jtag_uart:rst_n, spi:reset_n, sysid:reset_n, test_pattern_st_gen:reset_n, timer:reset_n]

begin

	debug_st_sink_0 : component Debug_ST_Sink
		port map (
			ST_sink_connection_data          => avalon_st_adapter_001_out_0_data,          -- ST_sink_connection.data
			ST_sink_connection_endofpacket   => avalon_st_adapter_001_out_0_endofpacket,   --                   .endofpacket
			ST_sink_connection_startofpacket => avalon_st_adapter_001_out_0_startofpacket, --                   .startofpacket
			clk                              => mclk_i_clk                                 --                clk.clk
		);

	cpu_v2 : component WiPhase_top_level_cpu_v2
		port map (
			clk                                 => mclk_i_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,             --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                   --                          .reset_req
			d_address                           => cpu_v2_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_v2_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_v2_data_master_read,                              --                          .read
			d_readdata                          => cpu_v2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_v2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_v2_data_master_write,                             --                          .write
			d_writedata                         => cpu_v2_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_v2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_v2_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_v2_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_v2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_v2_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_v2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                 --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_v2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_v2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_v2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_v2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_v2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_v2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_v2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_v2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                  -- custom_instruction_master.readra
		);

	eth : component WiPhase_top_level_eth
		port map (
			clk           => mclk_i_clk,                                     -- control_port_clock_connection.clk
			reset         => rst_controller_reset_out_reset,                 --              reset_connection.reset
			reg_addr      => mm_interconnect_0_eth_control_port_address,     --                  control_port.address
			reg_data_out  => mm_interconnect_0_eth_control_port_readdata,    --                              .readdata
			reg_rd        => mm_interconnect_0_eth_control_port_read,        --                              .read
			reg_data_in   => mm_interconnect_0_eth_control_port_writedata,   --                              .writedata
			reg_wr        => mm_interconnect_0_eth_control_port_write,       --                              .write
			reg_busy      => mm_interconnect_0_eth_control_port_waitrequest, --                              .waitrequest
			tx_clk        => rgmii_tx_clk_clk,                               --   pcs_mac_tx_clock_connection.clk
			rx_clk        => rgmii_rx_clk_clk,                               --   pcs_mac_rx_clock_connection.clk
			set_10        => mac_status_set_10,                              --         mac_status_connection.set_10
			set_1000      => mac_status_set_1000,                            --                              .set_1000
			eth_mode      => mac_status_eth_mode,                            --                              .eth_mode
			ena_10        => mac_status_ena_10,                              --                              .ena_10
			rgmii_in      => rgmii_connection_rgmii_in,                      --          mac_rgmii_connection.rgmii_in
			rgmii_out     => rgmii_connection_rgmii_out,                     --                              .rgmii_out
			rx_control    => rgmii_connection_rx_control,                    --                              .rx_control
			tx_control    => rgmii_connection_tx_control,                    --                              .tx_control
			ff_rx_clk     => mclk_i_clk,                                     --      receive_clock_connection.clk
			ff_tx_clk     => mclk_i_clk,                                     --     transmit_clock_connection.clk
			ff_rx_data    => eth_receive_data,                               --                       receive.data
			ff_rx_eop     => eth_receive_endofpacket,                        --                              .endofpacket
			rx_err        => eth_receive_error,                              --                              .error
			ff_rx_mod     => eth_receive_empty,                              --                              .empty
			ff_rx_rdy     => eth_receive_ready,                              --                              .ready
			ff_rx_sop     => eth_receive_startofpacket,                      --                              .startofpacket
			ff_rx_dval    => eth_receive_valid,                              --                              .valid
			ff_tx_data    => avalon_st_adapter_out_0_data,                   --                      transmit.data
			ff_tx_eop     => avalon_st_adapter_out_0_endofpacket,            --                              .endofpacket
			ff_tx_err     => avalon_st_adapter_out_0_error(0),               --                              .error
			ff_tx_mod     => avalon_st_adapter_out_0_empty,                  --                              .empty
			ff_tx_rdy     => avalon_st_adapter_out_0_ready,                  --                              .ready
			ff_tx_sop     => avalon_st_adapter_out_0_startofpacket,          --                              .startofpacket
			ff_tx_wren    => avalon_st_adapter_out_0_valid,                  --                              .valid
			mdc           => mac_mdio_connection_mdc,                        --           mac_mdio_connection.mdc
			mdio_in       => mac_mdio_connection_mdio_in,                    --                              .mdio_in
			mdio_out      => mac_mdio_connection_mdio_out,                   --                              .mdio_out
			mdio_oen      => mac_mdio_connection_mdio_oen,                   --                              .mdio_oen
			ff_tx_crc_fwd => mac_misc_connection_ff_tx_crc_fwd,              --           mac_misc_connection.ff_tx_crc_fwd
			ff_tx_septy   => mac_misc_connection_ff_tx_septy,                --                              .ff_tx_septy
			tx_ff_uflow   => mac_misc_connection_tx_ff_uflow,                --                              .tx_ff_uflow
			ff_tx_a_full  => mac_misc_connection_ff_tx_a_full,               --                              .ff_tx_a_full
			ff_tx_a_empty => mac_misc_connection_ff_tx_a_empty,              --                              .ff_tx_a_empty
			rx_err_stat   => mac_misc_connection_rx_err_stat,                --                              .rx_err_stat
			rx_frm_type   => mac_misc_connection_rx_frm_type,                --                              .rx_frm_type
			ff_rx_dsav    => mac_misc_connection_ff_rx_dsav,                 --                              .ff_rx_dsav
			ff_rx_a_full  => mac_misc_connection_ff_rx_a_full,               --                              .ff_rx_a_full
			ff_rx_a_empty => mac_misc_connection_ff_rx_a_empty               --                              .ff_rx_a_empty
		);

	jtag_uart : component WiPhase_top_level_jtag_uart
		port map (
			clk            => mclk_i_clk,                                                    --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	ram_onchip : component WiPhase_top_level_ram_onchip
		port map (
			clk        => mclk_i_clk,                                 --   clk1.clk
			address    => mm_interconnect_0_ram_onchip_s1_address,    --     s1.address
			clken      => mm_interconnect_0_ram_onchip_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_ram_onchip_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_ram_onchip_s1_write,      --       .write
			readdata   => mm_interconnect_0_ram_onchip_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_ram_onchip_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_ram_onchip_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,         --       .reset_req
			freeze     => '0'                                         -- (terminated)
		);

	sample_pll : component WiPhase_top_level_sample_pll
		port map (
			clk                => mclk_i_clk,                                       --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset,                   -- inclk_interface_reset.reset
			read               => mm_interconnect_0_sample_pll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_sample_pll_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_sample_pll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_sample_pll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_sample_pll_pll_slave_writedata, --                      .writedata
			inclk0             => pll_inclk_clk,                                    --                inclk0.clk
			c0                 => pll_out_clk,                                      --                    c0.clk
			areset             => sample_pll_areset_conduit_export,                 --        areset_conduit.export
			locked             => sample_pll_locked_conduit_export,                 --        locked_conduit.export
			scandone           => open,                                             --           (terminated)
			scandataout        => open,                                             --           (terminated)
			phasedone          => open,                                             --           (terminated)
			phasecounterselect => "0000",                                           --           (terminated)
			phaseupdown        => '0',                                              --           (terminated)
			phasestep          => '0',                                              --           (terminated)
			scanclk            => '0',                                              --           (terminated)
			scanclkena         => '0',                                              --           (terminated)
			scandata           => '0',                                              --           (terminated)
			configupdate       => '0'                                               --           (terminated)
		);

	spi : component WiPhase_top_level_spi
		port map (
			clk           => mclk_i_clk,                                             --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,               --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver0_irq,                               --              irq.irq
			MISO          => spi_signals_o_MISO,                                     --         external.export
			MOSI          => spi_signals_o_MOSI,                                     --                 .export
			SCLK          => spi_signals_o_SCLK,                                     --                 .export
			SS_n          => spi_signals_o_SS_n                                      --                 .export
		);

	sysid : component WiPhase_top_level_sysid
		port map (
			clock    => mclk_i_clk,                                       --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	test_pattern_st_gen : component WiPhase_top_level_test_pattern_st_gen
		port map (
			clk                 => mclk_i_clk,                                                --     clk.clk
			reset_n             => rst_controller_reset_out_reset_ports_inv,                  --   reset.reset_n
			csr_address         => mm_interconnect_0_test_pattern_st_gen_csr_address,         --     csr.address
			csr_writedata       => mm_interconnect_0_test_pattern_st_gen_csr_writedata,       --        .writedata
			csr_readdata        => mm_interconnect_0_test_pattern_st_gen_csr_readdata,        --        .readdata
			csr_read            => mm_interconnect_0_test_pattern_st_gen_csr_read,            --        .read
			csr_write           => mm_interconnect_0_test_pattern_st_gen_csr_write,           --        .write
			csr_waitrequest     => mm_interconnect_0_test_pattern_st_gen_csr_waitrequest,     --        .waitrequest
			command_address     => mm_interconnect_0_test_pattern_st_gen_command_address(0),  -- command.address
			command_writedata   => mm_interconnect_0_test_pattern_st_gen_command_writedata,   --        .writedata
			command_readdata    => mm_interconnect_0_test_pattern_st_gen_command_readdata,    --        .readdata
			command_read        => mm_interconnect_0_test_pattern_st_gen_command_read,        --        .read
			command_write       => mm_interconnect_0_test_pattern_st_gen_command_write,       --        .write
			command_waitrequest => mm_interconnect_0_test_pattern_st_gen_command_waitrequest, --        .waitrequest
			out_valid           => test_pattern_st_gen_out_valid,                             --     out.valid
			out_data            => test_pattern_st_gen_out_data,                              --        .data
			out_ready           => test_pattern_st_gen_out_ready,                             --        .ready
			out_startofpacket   => test_pattern_st_gen_out_startofpacket,                     --        .startofpacket
			out_endofpacket     => test_pattern_st_gen_out_endofpacket                        --        .endofpacket
		);

	timer : component WiPhase_top_level_timer
		port map (
			clk        => mclk_i_clk,                                 --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   -- reset.reset_n
			address    => mm_interconnect_0_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                    --   irq.irq
		);

	mm_interconnect_0 : component WiPhase_top_level_mm_interconnect_0
		port map (
			C10_Clk50M_clk_clk                       => mclk_i_clk,                                                --                     C10_Clk50M_clk.clk
			cpu_v2_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- cpu_v2_reset_reset_bridge_in_reset.reset
			cpu_v2_data_master_address               => cpu_v2_data_master_address,                                --                 cpu_v2_data_master.address
			cpu_v2_data_master_waitrequest           => cpu_v2_data_master_waitrequest,                            --                                   .waitrequest
			cpu_v2_data_master_byteenable            => cpu_v2_data_master_byteenable,                             --                                   .byteenable
			cpu_v2_data_master_read                  => cpu_v2_data_master_read,                                   --                                   .read
			cpu_v2_data_master_readdata              => cpu_v2_data_master_readdata,                               --                                   .readdata
			cpu_v2_data_master_write                 => cpu_v2_data_master_write,                                  --                                   .write
			cpu_v2_data_master_writedata             => cpu_v2_data_master_writedata,                              --                                   .writedata
			cpu_v2_data_master_debugaccess           => cpu_v2_data_master_debugaccess,                            --                                   .debugaccess
			cpu_v2_instruction_master_address        => cpu_v2_instruction_master_address,                         --          cpu_v2_instruction_master.address
			cpu_v2_instruction_master_waitrequest    => cpu_v2_instruction_master_waitrequest,                     --                                   .waitrequest
			cpu_v2_instruction_master_read           => cpu_v2_instruction_master_read,                            --                                   .read
			cpu_v2_instruction_master_readdata       => cpu_v2_instruction_master_readdata,                        --                                   .readdata
			cpu_v2_debug_mem_slave_address           => mm_interconnect_0_cpu_v2_debug_mem_slave_address,          --             cpu_v2_debug_mem_slave.address
			cpu_v2_debug_mem_slave_write             => mm_interconnect_0_cpu_v2_debug_mem_slave_write,            --                                   .write
			cpu_v2_debug_mem_slave_read              => mm_interconnect_0_cpu_v2_debug_mem_slave_read,             --                                   .read
			cpu_v2_debug_mem_slave_readdata          => mm_interconnect_0_cpu_v2_debug_mem_slave_readdata,         --                                   .readdata
			cpu_v2_debug_mem_slave_writedata         => mm_interconnect_0_cpu_v2_debug_mem_slave_writedata,        --                                   .writedata
			cpu_v2_debug_mem_slave_byteenable        => mm_interconnect_0_cpu_v2_debug_mem_slave_byteenable,       --                                   .byteenable
			cpu_v2_debug_mem_slave_waitrequest       => mm_interconnect_0_cpu_v2_debug_mem_slave_waitrequest,      --                                   .waitrequest
			cpu_v2_debug_mem_slave_debugaccess       => mm_interconnect_0_cpu_v2_debug_mem_slave_debugaccess,      --                                   .debugaccess
			eth_control_port_address                 => mm_interconnect_0_eth_control_port_address,                --                   eth_control_port.address
			eth_control_port_write                   => mm_interconnect_0_eth_control_port_write,                  --                                   .write
			eth_control_port_read                    => mm_interconnect_0_eth_control_port_read,                   --                                   .read
			eth_control_port_readdata                => mm_interconnect_0_eth_control_port_readdata,               --                                   .readdata
			eth_control_port_writedata               => mm_interconnect_0_eth_control_port_writedata,              --                                   .writedata
			eth_control_port_waitrequest             => mm_interconnect_0_eth_control_port_waitrequest,            --                                   .waitrequest
			jtag_uart_avalon_jtag_slave_address      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --        jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                   .write
			jtag_uart_avalon_jtag_slave_read         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                   .read
			jtag_uart_avalon_jtag_slave_readdata     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                   .readdata
			jtag_uart_avalon_jtag_slave_writedata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                   .writedata
			jtag_uart_avalon_jtag_slave_waitrequest  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                   .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                   .chipselect
			ram_onchip_s1_address                    => mm_interconnect_0_ram_onchip_s1_address,                   --                      ram_onchip_s1.address
			ram_onchip_s1_write                      => mm_interconnect_0_ram_onchip_s1_write,                     --                                   .write
			ram_onchip_s1_readdata                   => mm_interconnect_0_ram_onchip_s1_readdata,                  --                                   .readdata
			ram_onchip_s1_writedata                  => mm_interconnect_0_ram_onchip_s1_writedata,                 --                                   .writedata
			ram_onchip_s1_byteenable                 => mm_interconnect_0_ram_onchip_s1_byteenable,                --                                   .byteenable
			ram_onchip_s1_chipselect                 => mm_interconnect_0_ram_onchip_s1_chipselect,                --                                   .chipselect
			ram_onchip_s1_clken                      => mm_interconnect_0_ram_onchip_s1_clken,                     --                                   .clken
			sample_pll_pll_slave_address             => mm_interconnect_0_sample_pll_pll_slave_address,            --               sample_pll_pll_slave.address
			sample_pll_pll_slave_write               => mm_interconnect_0_sample_pll_pll_slave_write,              --                                   .write
			sample_pll_pll_slave_read                => mm_interconnect_0_sample_pll_pll_slave_read,               --                                   .read
			sample_pll_pll_slave_readdata            => mm_interconnect_0_sample_pll_pll_slave_readdata,           --                                   .readdata
			sample_pll_pll_slave_writedata           => mm_interconnect_0_sample_pll_pll_slave_writedata,          --                                   .writedata
			spi_spi_control_port_address             => mm_interconnect_0_spi_spi_control_port_address,            --               spi_spi_control_port.address
			spi_spi_control_port_write               => mm_interconnect_0_spi_spi_control_port_write,              --                                   .write
			spi_spi_control_port_read                => mm_interconnect_0_spi_spi_control_port_read,               --                                   .read
			spi_spi_control_port_readdata            => mm_interconnect_0_spi_spi_control_port_readdata,           --                                   .readdata
			spi_spi_control_port_writedata           => mm_interconnect_0_spi_spi_control_port_writedata,          --                                   .writedata
			spi_spi_control_port_chipselect          => mm_interconnect_0_spi_spi_control_port_chipselect,         --                                   .chipselect
			sysid_control_slave_address              => mm_interconnect_0_sysid_control_slave_address,             --                sysid_control_slave.address
			sysid_control_slave_readdata             => mm_interconnect_0_sysid_control_slave_readdata,            --                                   .readdata
			test_pattern_st_gen_command_address      => mm_interconnect_0_test_pattern_st_gen_command_address,     --        test_pattern_st_gen_command.address
			test_pattern_st_gen_command_write        => mm_interconnect_0_test_pattern_st_gen_command_write,       --                                   .write
			test_pattern_st_gen_command_read         => mm_interconnect_0_test_pattern_st_gen_command_read,        --                                   .read
			test_pattern_st_gen_command_readdata     => mm_interconnect_0_test_pattern_st_gen_command_readdata,    --                                   .readdata
			test_pattern_st_gen_command_writedata    => mm_interconnect_0_test_pattern_st_gen_command_writedata,   --                                   .writedata
			test_pattern_st_gen_command_waitrequest  => mm_interconnect_0_test_pattern_st_gen_command_waitrequest, --                                   .waitrequest
			test_pattern_st_gen_csr_address          => mm_interconnect_0_test_pattern_st_gen_csr_address,         --            test_pattern_st_gen_csr.address
			test_pattern_st_gen_csr_write            => mm_interconnect_0_test_pattern_st_gen_csr_write,           --                                   .write
			test_pattern_st_gen_csr_read             => mm_interconnect_0_test_pattern_st_gen_csr_read,            --                                   .read
			test_pattern_st_gen_csr_readdata         => mm_interconnect_0_test_pattern_st_gen_csr_readdata,        --                                   .readdata
			test_pattern_st_gen_csr_writedata        => mm_interconnect_0_test_pattern_st_gen_csr_writedata,       --                                   .writedata
			test_pattern_st_gen_csr_waitrequest      => mm_interconnect_0_test_pattern_st_gen_csr_waitrequest,     --                                   .waitrequest
			timer_s1_address                         => mm_interconnect_0_timer_s1_address,                        --                           timer_s1.address
			timer_s1_write                           => mm_interconnect_0_timer_s1_write,                          --                                   .write
			timer_s1_readdata                        => mm_interconnect_0_timer_s1_readdata,                       --                                   .readdata
			timer_s1_writedata                       => mm_interconnect_0_timer_s1_writedata,                      --                                   .writedata
			timer_s1_chipselect                      => mm_interconnect_0_timer_s1_chipselect                      --                                   .chipselect
		);

	irq_mapper : component WiPhase_top_level_irq_mapper
		port map (
			clk           => mclk_i_clk,                     --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => cpu_v2_irq_irq                  --    sender.irq
		);

	avalon_st_adapter : component WiPhase_top_level_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 8,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 1,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => mclk_i_clk,                            -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,        -- in_rst_0.reset
			in_0_data           => test_pattern_st_gen_out_data,          --     in_0.data
			in_0_valid          => test_pattern_st_gen_out_valid,         --         .valid
			in_0_ready          => test_pattern_st_gen_out_ready,         --         .ready
			in_0_startofpacket  => test_pattern_st_gen_out_startofpacket, --         .startofpacket
			in_0_endofpacket    => test_pattern_st_gen_out_endofpacket,   --         .endofpacket
			out_0_data          => avalon_st_adapter_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_out_0_empty,         --         .empty
			out_0_error         => avalon_st_adapter_out_0_error          --         .error
		);

	avalon_st_adapter_001 : component WiPhase_top_level_avalon_st_adapter_001
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 6,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 2,
			outDataWidth    => 8,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 0,
			outUseReady     => 0,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => mclk_i_clk,                                -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,            -- in_rst_0.reset
			in_0_data           => eth_receive_data,                          --     in_0.data
			in_0_valid          => eth_receive_valid,                         --         .valid
			in_0_ready          => eth_receive_ready,                         --         .ready
			in_0_startofpacket  => eth_receive_startofpacket,                 --         .startofpacket
			in_0_endofpacket    => eth_receive_endofpacket,                   --         .endofpacket
			in_0_empty          => eth_receive_empty,                         --         .empty
			in_0_error          => eth_receive_error,                         --         .error
			out_0_data          => avalon_st_adapter_001_out_0_data,          --    out_0.data
			out_0_startofpacket => avalon_st_adapter_001_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_001_out_0_endofpacket    --         .endofpacket
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => mclk_reset_reset_n_ports_inv,       -- reset_in0.reset
			clk            => mclk_i_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mclk_reset_reset_n_ports_inv <= not mclk_reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_timer_s1_write_ports_inv <= not mm_interconnect_0_timer_s1_write;

	mm_interconnect_0_spi_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_spi_control_port_read;

	mm_interconnect_0_spi_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of WiPhase_top_level
