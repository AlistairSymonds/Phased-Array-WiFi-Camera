��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O�Ä��/����f&4<LY�~R&i~�0�q��Y�~��<���Dp�Eñ�����N4�[G�8����og�=υ/�3E�D�0���?X��fQ j����*acR�^���WW�S�e�?�w)���[�a�y�R*��U���� �zzN��A���=iT]�8���@���`��\m*��̬��)��n���٣���>�&oԂ8a�L(Gy�F��3U۹FX�Nv�Ѷ)_�e�����lU�՘g�FY/��T�s���b�9ܧx/P�H�l6� ���r�C{[��%y�Ab�=�s 2V9�p�P�"���/6�E��ɐO:g9k�x'��wv㱏6�	��euW��)@�V���)o��T5z����%�߬QގVKѥKb�a�w�����I�Gk@S(�X�̡����Q�3+[�rt`�Р�@J���']����C8��A68��T(M7�ڬC���Nu`��2
�pdߖ�o<(w�詌��)l�k�߻l�x��J" tJZ���IT��]_�-�<Ђ��@����.��rW���/��d�ߕ�T�vK2�;���1}��Y��)��f���I-�蹞B4cN�#~��,���om�h�;~ů7���DLɅ�4)�2�Y��i% ��"u�o�C��A�NM��A���b��#��"1
�2��a�!���8Ko�I�	-0��̈́����X��I�x�T` �P�^Sc)c���g�(MХ�\!p<�2Wk�P8�V�̸/�v��(�C�o
K�R��v`���7�f��e$4�BU�D{���;oJ�V��J<I����7��8+V�Oj�~`�nI*�E��v��M�zM`nN���
#�k$��͖+{#S����#Z�b�|�|3��[	B���Au�[��^�Ѫ
!/2��XM�:f^�I���߲4�f�=�bU'��M!<�(z�V��N�v���o�	���u�I�0j���f��(�O���7�6�@����'�&�'v.�������ئti��e>˛뚖=��k�B��)�~������Oe #
A#%�<dW�f���.�	�z��U�e!p\ Ķ��G���Xj�b�q	Ce���R�dV��8:#�_�_!�ھ�X��Y!�ܪ�_�����17zN���p�I�`�Ovs��b���:5~�q�0j�\K��BD3�{I#ěcB��)��� x���`���Ʀ��Y9��$�	s�P��!z����ݛv��KO�XGa�ShL+�����X�8��g;��L�r�v�]�a�P���X6���<߫J��zo}�:�M�����8��e�}n�~�k[������6 ����{��@��P)���2��2vK�L:V��X	�RA~���.rIʀ)��3@[�{���c�ٿ9M���t���iO  �D�2e�-b���ޚ����#�Kh$3�G�W�$:�T�t%�_ѐ�?�{y�O�dr���E�[^C3y6�	���v7��=�|����nE�b�ԇ�vONh5O������J&��<�~�T�m���Ԛ�I��瑊ߙ.ظX�:5�{1�J[��������9��V���ZwX�s���.�� ߂~1�O@Ű2@		���8
yM��q���^8t^�Cf� �}�6b5�$y.U������L�r�����y�tJ�l$�\4��z�޲1�%��m��)�.�я�6X����
������p( ���y��ܸ{6��m�� r���d��XWэ�����5}������)�'3L6ô�xhV)�R�#�/c[-���<���-\]�����Ny�@�M�Z�s�C7|��Ŝ�_%�w�%9�ݮU5=s%oVv��)�����s�09:X��4�m�,'�%6}c�����d\|�C�*�7Ϊ�&����zs�; ��7��kl.�?�������*j�ϕ���%��R8��*�0�}`<M2���w��4E"AC���r��`��q�E�NP���@�< Z�a�v�|�C�WxN�4��\j��?V�y��L�Z�l]����&K�f�1��j�qX9&i�]*�knDu=�x�9����r(P\S=�Ioږ3�@���'�ó��!�XAv�����(`�e\������&�k�6���� k9G�V�N-�9p��|�{�☾�_"����,>S2�h�H�"#�Y��e�
));E��
\��_ ��q|���Ҕ�1:?��VFk��#o��?�⷟m��o}���=̷��A�1'�(���6LF���Xtb��º� ���LBfl�쵫%_���zo�9��-���S]������Y�t��}�MFp��-�?���r���tV? ��
3�,�w���	���p[S�7ì�E�5�f*homC��s'�~�5���1�b,C�m$إ��N����b4o�U&�^���\�D@�r���/5�Kҩ(4�z�to+<���ZP:��?� \lh:��(�?��I�����@������d�PU��1�q睗���*nq�O4 ���{���x>(b�m;�Xo�EG�t��@�b�oj�wiQ8�-�Ș�n`��S�T�����2_�_�c�pS�9)���I��(^�&c��w��.	�M{�ˎ?��!���&������L�e�d���Y��� `dS+8��y�;"f^��F`�V;�V��w�U<�@��c��?�Iٴ�KY\[na�M`7�YkoKnw���,��v9��g�������!���͆�+?�h��3���v���y�`TB	��:�g1!V���?b��L8;�KS�m@�a�<���\�����^�u�6��\���J�!�� �}�02,������E
���jV�!�"E9�8�dRc9��t�,)Mڔ��E���-�I��$���s���H+�y��m���.�1��n-[d�˩3���s�>�-�Q#�}��Gm/po)��˾� �M]��/ؤ�v�|u��ȳ��Q�VZ��w+��I�2�q��,�Y����ȤH�;t)����
h��V3��~��p� ���V �  d��U���KmS]O�c]�qNO����)"Q��Ybj
YC�#�Z~Aɪ����:�o  ���SM��R�S�6x˭匛��q�N�L��;
�L�6l�c����=�@fX�����S+pG����J]Ux�4�$�6�G����ܸ�	�K���X��\�s��m脥��&���Qd*�R+I�Lw6���%�5y{W4	}Z��&�6�6#�ہ��
�w�K?u+>��1ːّ$c���D�?2N_�����C^�:�*FK��T@���~!��Р<��I���&��,٦�=��@,ޢ��µ��m!
su-�@�%�(�('N������ډ���&�q=KP~NB�\2O��t	���
,ҋhM#��.Jl=�֤�b�r���_�R;H�3���vl>컊���+5�Y�	y?Ο	5K���MԘ-�<p�ٯ����/�x�8�y�rg/��
	�;v���G�b���#cF�l��p�����b�}v�$b�$�^��V���Ԁ��lc�e #���x�,�y@�ˡEE�6��o�4�L���I����7�����v�ﮡGM��9Xs��%߅���I�;�����Hd��d�x�d>�����N�"��f�U�K6�d�;�9�_��W Д�d�ݞx�cc�8PKfC���b���K6Tta'{Nߐ78�V����|�X���1�{��^�����E��@��9�Z���X�1�N�T����T^�?zb���+(96��nN(�8KAk;��,�@P���Ę�"��~.,�x��M�����D���S{c�X�}� ���Pz�˾��e�!�B���V�h�N��Z]R�5����i�� �LN,p�ö\
Ң>��)���-,�vTn�\a����p93�4���v7dj�%�n2�\��9���q��]T����·���n����c�Ӄ�+����:��3���g�' �6A竦��:������]�m���ro�<����j�+����K� A�CT��SF�6��hƏ��)@�y�q>UZU�䄏�ЫA��~_�$�9�'�^&��Zp��R�Z�=�Ņ�q�L�`�x7��te�v�C��D(�f�-�d����r����jEJ1D^4(��aLX*�Ł
��u�ֲ���x���֐�&�&�d�IS��L��	