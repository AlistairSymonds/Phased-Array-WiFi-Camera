// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:25:54 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Dui2uZyVlgljpvCUmFfg4WU6eiPp/R3c3ZMqYl3V5G1HHwRnbF3dHkjtDNi44OtK
39rlpAmC/3Q9C2dGDkUa/AUtLH53w5OPpsY196jluvtlT5dEGW81MkkglAj5rcMp
RuFMLH+1zvr6wVBlrwmWRzORmIDPHRQexh50usv9XT0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
P7agOSwFPZfhRttxZ0O3HiGnJZC89lqjCrQN5fJxvNf6nCfdGmKx+gn/YD1fFrD1
dzUq6isbwO4wqcPnO0O6JooTcCdoMVslstka/uhhDZp9RkGmbr/3dIRZBVRHMvtr
RkbBT3iImx5pQBZykuESac8Z0AgGAxIadEbugWpSYCOE0GjtSzBwfCMG8rw+L+Ar
1ISEabMLohLXbyLSWgeblWHKDYfVzP8nqi1OyGOFGz2QwOiBfxrEeOuP/D0rbNxV
AkAHpTRMXOL0h/LbGyEDeC8jY5i6ZmqD4ksdLWAR8cNyH9C/qMBRW1Th5vHLrhmg
3fnErI7sOuIx1uQ3tNtEds3qV8/0chMM81y8RxPCb+mUbqQ48Ma1zyzCB1Xf1wjC
kwbOmXMXPlM2TR+UvwBqyzCuXZmSR5rxvbM9icDwurhBWbogDcQLWmR+AjfDUYfF
1y3GDXWw+05WIJujLZHk6dgFQms9yVG3qbvxBOvIdc91CVzrwv+shujEfYEEexz6
aJXLLGwWpiCBsb46/aTliKJC/7zJ+drpWAa72HRom8BN5ZLQMUOCFw4fg57YMm10
OwPRAyyz7A2XMrGUDxPIVCFZE29cvcSoKkA3R+Ujxaws62IS8xTBHCuz3RDQY/Fd
4FsrnW4ZLJ/Zmk8RjaEWhYMhqUFAhkdXYwEJeyeINb9L81ZDwclPJwvPX56A2+oI
OqlEastQWjg6HIRMjFus7K3fEqaTeaA7+4k0GXIW26gTMTXyM0DJ3cBNkaTVW0Fu
RMSK9EPuvDK467vcX4B28Ll9QdZGshhOhYaE+E266sAADE3dGXyzjOm86DPXG+4x
71xwwPBs7CfNxVpyMeDwXDWYIeFR/mADHNq1BZUuqFtmvIIe2R4Bj7xVXcIQ8dvP
+SHGb0b2Aq6aSuv8MkOGxGjA1rZR+DRi6pFMTWdqoaJiq6LaL9eO5CLwrkdNljs4
ApqAawYQPClkSvFBbo31p48Oc4LaqmwDAM/it46wSeMjE6+7Dbdg79Fl+xxMHR5z
P1iQb4lhIDVj+pZ5NKEBBFPN+q+rc1UhgT7ArSqVo8urQpmAMhDKJV5hGgwl4zGo
UCzn1ED1EfGtunZpW/QOnVj13xiCmKPRF6L2gdNZinIQz6UGEDBYLbCKJuMDYn/R
CQSXugmBTMMzOml5HnLrxlqonaOJuf/tmXq1aEMnPnt3yc8qYjI7f0+kk059Gx05
J8u7zWi7fSsvZ+Ik1uLfyFKUbwE+tHwlzw3P7rywXUpjb5nV5pKllufiom5Njnbl
X3jqM8HWqGyvKIy85HR7sHfv1UZbJCMiqAigiUuCbySyIbLW4n5DqrTDNTVxTj79
AxnTymRnQoNbKnTRrusJs7AEe86lfwasgbgpJ8AElyOvNSDfc0/h56jIwoIBCT0E
5rL6feiwegLrNsrhFIztaXODq+chZaMeDVkq+lNqkOnAePplVacO/BVAYB2l10Lz
N3O2R2eFSkMC7bj1izhvLRS0JufaB+1ZVGi1iEhA4QAgoQX7PJQnEPYq/syv2zMV
Hhl0UuiujBvsBpRIkB/NJjk/SRr+DmSzFBNbyEHhY4lP5gn5EfzmAFbg47BDQ6MI
NjNKdYCc5/ko1mQxRplehMnu8TBhbDq8LMVppMW8RFyVFp6OiP7Wuwx6dF4z2Aqw
MlKjvdzyWpleHim5mfxpr148/qjwfVMizc0OaE7PtiqCeA1wpNJAZLHYiNFIRO+S
1Dp3xVzWgnlC5jiQlqvLTbMyTqW8DJNOYLyaTT+hULg17OOuEFXiW0tI6Jwb4V9L
Q8L4IxzFi9SBylKmt0ExDXfoQx1g9NQ97s/incgzK5YUHoFQhwQbJtmsYjsgiTmj
bs+Yk6vVMa26yWNQ93yWWcAhlhk2JT64q8BufwVlWjB4v2hswg+gcbcztMKrWCKv
FfwhM+rqhu5lYaVwFAU4ywOTW/aSyhex+OlflpDONwsJ1xQmODQ4UgpdDtpy9sWU
hB3v6YkXgpyl51icP4lig6/JqoEZthqEvGBivDdfzfFnOX/jKpvKFg//Ax0LgFvl
oTzf2d3JF/dsR8GFUuvDTU3dM94zXhrGnF72eM3nnwBVsfhEnaBt1o7JLhd+C0bW
1eT76b3w80NqXudBbt0Wz+Pt36BWtOZAxpOQ1iVM0G74/QripXLDhH5x66Eqbyjw
jBp+Q03UNz805t6SicQ/bq57dHAllmgsBwKc0l2J547zizHmIG9/J+2OSf5BPb0D
owqrS8jJzEUY8n8z5y7X6Bm9JGoe23y/YnBrCu24gfA0WXyS7dTeBvX7x2yR22Xm
c37VnHDff1EGV3S/rlK5Q++aZa8S5My4WZMHj5GY4kHAfaaFhSdScQYvZtQwiqrv
auMh7ZOnHtmhgSHO9xWoTuFFqpoJzhUbkWzPMOxbIwIamlB6B9SzikBNa+05Fz8n
Qve7M0MEoVAbJeHZg6Dsm/HnDjcWTOXadsht/8fhz+C+2JyanYSX09Str2f/i9Jz
cCjXNa50HfGZCWr0iw0/z+D+NTgm3+sTUsOB8f2iz4IfXKsTxVdpOt1aQx7IrA8F
eG8t/jElkB2MtIPza4qmwPJX2gz2fxhfzV3gseSNn/iez+Q//hrnicTIjyDdITum
d2r8uAqx92k86kesF7TLiHu4giGVVBTeUrULEG6LdJH7qxt+I8k4b6G+NsGakxiM
DdyaOGqVbBIB/deT+KksBPxFcuN48UrdAJhFKA5VskRDhphlqHcjnVghxX8alkad
YoB7r1v6+kt+PlsIRRQcw6fNm90JBRc03XaKrIyfpgMfS2Lg/OM95ROwCg8MMI2p
N8P/yWMXqNeb4AzScbeFplFsZmGIYwrZRm+JO8N5BMep4pVuofL3HOxJADUkfMAc
Y1iQohJ/1bMgRHt2Whxv1k/uiJqP9I1Wqp2gyd8fwTzo/e9FYoXTxoqZ7yD3mQYo
22VMYItszCs4EtErNqm4Qm3bZw1ikm2b7JS63TPXYivvdunkpoL2jyGZpXVwXGKF
8iR4t1nTC0mBtRiHNCxigBxy2QE8a7AMb96tqeJhGgyipKUlPTmnfXGuBlSS+x4h
Dzqs1rGRFnMKWOdMEVflfwOu5WP+Mvsa/woMU23OaV1OiBbjbtHubyQwchjQnJRU
nE4BOQ9f1DhC9brU33OEEtVPQHGmKO4aVXs6ysWi/VIibqxFWNlMt4uaUzw1lGeV
UGk33FYmzWgGqLE27aX5WnoAt+MIlRpiwIr4mCuuxQ2vz7Eb8qJhbNjv8fQmRJYP
9ofztZ1d+RuWP/raL72eBpig/dluatDZwJHusxgUPkYWYdub/iRLqXirf7aAbIct
N/qF9/MIigJ/jyir9EuV8FTx1HQViljJcYKh2OLTF7EkpNA/JjqtFzYjwectGHQZ
BPYNpcQI5Yvv4/c2XqtvgIfNsy5ew/8/I+7/E7F7k2G3F+s3rdjQgtiQQ1lcFPtt
elenGfKNVkfP2rGZtgN1x8SI3gOtX1BwdFHMP+l7Y2TEl8UxbnTxdPJwvYzUnwAz
y5Q9cJT1dMJImCXFrjZY1X+SRPfjVC5b/MY7SwA4rGpaD6Flt/iQ9p+FGmt0jCqQ
0zpA/llQNWHsx98yMmrbjhOvi5bo16MdBnhXqFRDh0hGMk2nOZBYRekRSUWxCvAM
Xns2M5t6wMsQqaQ2hocl7gYAL97ORejQ8/tq5G6GdbY0ntnJwpBBkjN42onUYcmm
nu3/Q9FHw9ptYr94SS7JZNPdVI5zHJaCbPS3q9YOzCCqyN7/NMihJteeWAEvEL2s
us961p4MZHuJDU/yiGS2alJmAhUOama+og0tMSoXtTwDDolltT/0CHaDAU2RtsQm
h8G4HRJoWbxbVmS66gTLBVidRmBUkcwIUKRtuK59Nvmmdj1sOc0q82oodW8wIlyd
kmtv+KFBEvgm7w5P4SI9njtzL5aHXjL3yJP9pFTzZojrXXShigek1q/lLuICJL74
s06l6m8uJGjyvtoO5Ec9fDguqeedXbgKOE1rH3FK07Hksf5pIevnx93ySdA1JQ/w
cvG8R7B4hr3D5U5OTYutwAImnN52r/PejWLBJ6BIXlYPTEFAq5nxdy3MrJ7x8Jaq
Nk9+a5E7S7fgQGCV+dAQi13P6rNqs11EiyMkLpqNfoxBeLJxOba4+TvFtHzRIuDM
MNwSTofNE5YaGCD7787nC4Bd1Fhrssr+S9B+SQUsflO1Rakzo5bdqopxHDQcGtT1
U39G5uPen4tqovU4/Gn4cb9dVLl1FDrXjwsy6R1fK0qXUeXZIPQX+SZT+d1C+I14
kgQL6DLQ28KyrEAvTTX72fHThWxHOljen2J7hSJUDL939uz6ADdHKkJWLIIXK5fs
1cwY7B0oNHyzF5NqHETqDgK0XHWGi22aP7nmPq0YdY0cxx4EjHU+QnFhpxrux5tj
/A0Ni1k/ulPQUWigUGfeDoncm3s8UGOZRN7iirtcnShZvbxKp1EVS5I+UMnAnshb
6KYCUXtkr+gMy4Z9ZkDEKKTvqhp0rfM0MuJKwav8oBMOIaMDdY9hzAlnptpPrfiT
I7IbXTsU4L/IOms5YQ00Eamio58tlQK+5lnUfbeIAJi6UkjuCdtuUBo0KnN/taTO
AAA1TXeBOphZ7PdHU6QB8dxec0bXIOWQhG1s76rxdDK57s1HrEIEkYEkylhuNuYQ
wFuRDE7jwi3wpQCAQ/EjrO78J6D3aWb7eyMRhSoli4c9ROpn7oGSmsj7bS3IcAiU
iuv/lFIJVJq2I0MM+007YNOxocMM4H8bvCY2N7tHx6PaBkkWJla3uNrrsv7tO+7R
QWuJNWRNIFrDV2QtfOBc3UmeLCV5XSxDYeJONE7e/SOu4U5wyOWo/5pzjzrMSmYr
6wdBkxLHkwnup0AB9YOgwDKnzdUl3gTz+p9YGiZE/42avxSk7RgfRdcLr4JjnNAg
d1vuow7bHva5HFRc0DpI+kVDYlmqFOxKd0V0Kjh8Qal+KQCgtZV7b9Kq4WR7enu2
Zi11aVAMgyLTKVHw4vqEOfSoO4jKzGQHIyGXkTUf4dFtKgEuqJS8CqvY1cqniBwR
ZHfDpGK35D6uGK9TD/tEL23rFFe3ykKBw1PUiKavD8KHGJgMUROfp6bP66CfKgtR
y67KE0iO+ECoeBeEQtJTkw78XeFlKCYROUaF/0yBN2VNSrn7Jf/tlnFiAh1+KA4z
Y/TBBOmC2WM9Db393n9yyXpd/fB18BzEX/4MtVhU2vHsz0FFB/WGomdP4MkjtYhh
a01eB4wBKZpZgtTFweQ9/+PAcht1YqUbG+i1s8JTyZXxVm5FzGu6GX/LFIohODiy
+Lrhc84iYBBpkF+n6S3sFO7whpxsxcJ+3FyzpEGV+eWaHwU2SlPL+3pFlq+8unIx
irss3PDVSnRqM8lbRve/yp89wYrQXXQW7E39hDBbHlHuHOhhNJUGOJmF/sywVBev
dSLBTlr6Sxs4VGcecw4R1eM8LvYyNIEP+I+xuqF185vvCWhCiD6X57UaYR46CYK1
7OB34BXQ0OVLNrobxQOoBgsQowQOjp95qYbo2s9vGeV8X9PlHVL/og8oOqNTocDM
wwHhI2wF7nzCYfP3054W9Gmn5NR1nbSO+NxCIb1pwdA0QOjVXFUSSh+zj+C/S2iP
hKeWEJmd5ITm/f3aE1ayshbqK84WcmStrP23ziMatk8+4UbVkfpVUDl7nPdUDEQx
DhOfBQn3B0vIIM7VC5sdd3sXqh/x+fS6itNwxDeyHfDQHjk8hsf6C16RzVHUAkzc
/81C2IJdRlhjlT076GuOkkPDJ5ooIHQ8EPbdPFYvdNVsSmF0cHng7jCpFfPT/iv5
k3wpwuvXNVIm6M39cfAlJpNs9ijlsKALa9rp+u7vW3b4xDWs4FfoAJin5uqyAYRA
I+221DMIx99FuOBfQdfZ0ReD5fAN9ufhU+ZUmKN+Ma9uWJt/4YXL+SJJVnw2jXM6
XcEyCiqr3AEQXZAt42L30qkZ8802ioSMiIyUxbHd+ZO8KGM90aK2l46UnDIDZOX9
q0LT2oCjkTM6mad+hTJj+muM3NmiDHE0U3FqEd3C0Jh9G2b0r+hvg+7Tn8JgzjIj
+trpNYRGCp7pvoAKUHUpGD7fncKJm8otYLvF1AmNONN/Cx/U4NJ0W4lJECmXIqkG
gNCfPoZHEc8FpR9xYYailubmia0K70MyfS1Il5aubu1MwwcUAXyV/y7ug9r9+pYa
mcB67PWEOONGj5bJXi0gjLUOA8vHCbkZEJYcbFuAQLXM56jXpspFNioIYTt9teZ8
ygcX3URbpFDYzF1cXFAQEgIDZb2pdGeXKYMg+8RIYp5C3VLW7tWi39eEesvO3Bem
X3+WuEqt62R3cCcMFTwCzqTZzmcwA1/NRvJsNjMq3Syf0adg4JQeiWhYrNFjm3ei
hItUgC66q5XfMXQAKtkNORbexh6lymYJcqmAo1p320jl9QYpAolLv0zu+6dET5R9
druCEcQ9yiJ3n5Ctfs1n2zQYaGUtXM5YLO1v9IMYP7TlfWLh7omdADqwYQEYIsNj
INMKZ7MkRMcL3e4o0RcWLmitnlCGPQGC5KT4A2rjVxCj8Wh9k+a8VsYAqpVCMAus
bRUeCv1Clq8CmnzNdGnPBhop2D4Ckon/oXW3LT4L9wTLFwWCv3AnHJuR114yxdsM
2GywrwDu6iOCHDNdJxYlVlGqMET4MWzD4utu0nX/3EejwZRBOL9Ib0IvpZ44ZZnm
MVPKnMcRnOme89Pmk03ODEuFFsD4bByfHVounTs0I0NE8MAWMUxUVENf7ZVWkZK6
LR7ND+m+9NuApfcBspXSonUd7guz01XZ+TmuMXLnoVfEGBsxEmEPW462wC4AkqdO
VhYUnJf4mc9aKRUi+4B26Ixs3pHM+YJEq/ti85diVxyGMCGtkGaWfR2tOvKYpQWx
Yb3iA/NmpRSPrxFKsZWuKtkyqFpA5s6umm9sRO6zaVI8pp0Eh+2SWDR6EUHakNNU
N7Q4q9eSkoEZAWFpMFKdvpP0GxcXdThMjkC5Dm/R+PT6BfItZEI9wjItHbS6nuDK
mV3A0rA0eAW7G0NMmC8X+qOxe3tjSeWR48vwoA7ZvRfEwJ/+/DnXgabu9ZyEYDAj
myLJ1sbULqtk4LelRc8WON0uWHjrrEqEOKb8k2mxcwLf6FAzfaBDQCqubRhbTl2g
Sny6Qxi7XZURCacNJqkjB4Ps9BmyM4B+jRK8VIIF9Bf27f6rpeJ3IY4yYzqsIGzu
CezT22qNVEd/3+BQFQx750QlqIG6u1vC4bchxOrg3leSLvAwZF2wGqh2mwN0lsCx
LIzeypDPL6dKaWIFCn39ydARUl3W2oOG8R1EY22GGffJ/GYlelyKpqUMkogLyCQx
EMnzxKEC6ero3PyBWubPsBRAPxqFYVlAC5YFMR0Of3C76jBhNL4E0CF7SJ6E7nsz
pol/+lpJ49yX8Mv5TIhLWtA+9sCMaExgxhGm/1+hi0BEvZCtbTKEhKb0t8S3YI/d
XEyE0ASMCYtWTT8nlDfHrkvMHSm/a2nvrh8zmzqWaQSSPNEud2ZAb+vpY+3Ru0K2
dkH6JuHeAAJCNcxgzU4WVVaIvQvkbrIrzTy2kXp5V8zk2sQ37DJoDac8xgPRf330
Ip7jYwbfw5zmbfO44Kj+eo5vh4DPM5Sz21Ez5DuowzEqrblgV4OiK9yqj18WcMbR
zu3Q09k0ufxHrTsX0MwIC7PVtQJ+LmOFe0GxknUpXbcukpnHGA2B6hMljQ9oIh2e
G0XYwnZoC1HL6QenPaYGzbHo7qSOhwx5qB7qcf8mCvQ=
`pragma protect end_protected
