// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ZgWTrgDPI7z10uCyOs7VvB8sXv/8r2+zB37/dkRr1/wnSzA8HWvl5KRWJych8N+yXKRNZ13K8sfd
jc/Oo1UkK47kXVHv0RcMb3Sm1OJpDcnQwOets396F/qvMJ2v2tvsJW6ZA6fLZQBH8dVUxURfh/Kg
SrFrJtIGEjEyhtmwJNTDZgosYaFJCahrBejjLA/99sSr3HQ41zt8YBk8b66CvEQQlPZbmzR4zztD
HV02nKuX2sf9CByWo/sSJaDxefiNw4E2/WTlIlrz/5Dwns4NZ+UxaRuM/PFpSKrQR4RcwSu5qYrh
/e4EGVw408xQ5z5VxYr7knzDGV05PqXISOicRg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5264)
ZxSc4ZMSyNmdcJGcTOfU1cdD3OIa9/G+/0Jj2om4VwKRjPduOQCbl9OvkiADB7/Y1zF1DBFi1lEk
hWaVJ0OhiAeqMgpu9HtEhYb9mapgvK9wmsqZq8mtzOzB0BIaVhmG7C0Qifk9T5Cgp9UHG7SkOXde
Ex/fR5xXXb1zyFOQUqXfW/F8zURkqR/9KAaJeHl0ivx7iadsatAkIFJagQn++Xw2aShMQhwlmBbY
rAQRQJg4MNDjxvMS79HKQLIfwuz+KUqrJUi5ckmsGmmSrf5+1NoZQqKQsZRqNsDaUx09irXiXZy7
U/snu/eX5jbifx/266NLOsvJVclJAOLDeI3erNLdD3Y3skUzlHQ7Uh5WMFpZzHodY6hEfDNpixc0
kr53qgwycpqd1WorLvIIVTolbFgtzAsunj9kLzefpsczwhC5eSaiq4+g/I8aJckHpu4nR2GhCFde
Hl42FR6HCszwhLjiQOfsyiJOloYEtyZnHFfRVPBTd++Yf9XsLgaXBR5hJMPI5YJENITDd50obxeg
M90Fc0LF5+PxeJg5fzVBMJ8Y0bstw6JwIRM3tYJOAtorIOM+KthnNKCrEYjRMkMusSM/9Oe1IzCX
RWqrSr5q3c+YPbpK2V74ooQg/mTcBE/CmGxM1GqKow1NPD3Wuk5IWFrX3zHc0SxF36CdadXlNtrM
C6X82Z6XdekKd3KtyvxC7UpDqjHwS4SyXoDWLhnCjxJK7P+lqB8yzSAxeYVp0MGLvL5PX01Giha8
tsZIC58KG6Di8a/5cWWQ3lXjLFb4VrHU1OP/ror8GchNru7Kl+MQaeP2AxDiAwqt44nmpB1KudTj
qMITBnD2wE9+wLITeQMx5IY6RfbbPf0z9NjKO7LFr9TxU/11xtfENFGNnx2JZ9uwoIrP3snah+hy
XojTiPewoskvvbQ/3uyXe3FofFN4LhJ3xkrXGPd13tODTfLsVYzng7dbLvKXCVUEs0eI1umFOVb0
apHFLwcCMxOU+oh0wEWQ+0v01N92YU+5hY4PxYbuW8SAodhVvjLawDvK/HaOe0MPdC9r4MR/zdXi
hBAx80YKR6aNSpEcIZ1zkz8xyB1Z+ABEWHswyNqDScxiZm+CDORrXZ4raqn5aSvhVzE5kHaKsJni
yooteZkNCG9YQIfaCaLdAAs5zlr2Cyhxh6FkHMzsW0RCfbDVlFnXPMWR4Jn2PVfY4D+MvnXIjOkT
ZmEVoeUqZ6J2zz0xGsI8EL7iwfRfdVNEQX4jJZEcgPunXvwrDEOmsdVu+U7rFGtsZSz6n0FKco5A
33zd/344HBWcJTbhjBKJaiU06TCV5ErwXmMzW/c3LiY+Y4N4mNo8CrhY6yZ5eYRz/iyTTKqUPJ7V
2MaEFzAKRN82uiY+ZEtiomnIlErhwfdKR6a1fTGVzizlWdAo6GxjB6N6SB1W0m0HuRI0TAsLisw2
q1IeJ97cBMy0Pl6kHSgX5Vl+QrmapQAod2WuzbMRfXK9PrQPWoSeFWl+Bi7lvKsYZ4Frep8+M4PR
ruz7+Oy7bwtE//n+1HJqpzk92sWSHqRnLDEBv7mNHMu9/YwO1tL6dsPCFXyxi8MognVfUn90f6km
j/glizzat15DDec0uNMrNaTg3LSO/Xcy7Mf8gMzrpGEDF/O1hOzaC/nojKbXVPY5u/yrf6IASbPR
UI80UFBFF9oP70kMGAENWSPiX7FWCFBq8Cz6vdZOFhsljf2R+AFE3IkctRyAJjbNvQNuQ+2yB1tH
ClpDrBHx7gNZ8eMnGH0H0LKZLgzlqNR1bsSpzL0nYqdcWTvilUC/Q5z1vCnblGrjpp50bPqXV25N
hpLJvUOKMkKikYXiNFQT2tf43GEgGVPD7ByURlYitGH7qLZYAmN00rhmAU6eY5azji3zE9KJaHrr
QkZDrGLxdbHhQLN7HnFIyLakedtulroD2yF0SCpvifYNJrFV8ZMlrRsB5et5eCtC4s4zmZ8n018O
dHkvhb8Tho3PTd/3QayHOzZdDdoPH8ntX4aULfPjN3WpJbvWweenuYai+PpS+MIQuPTB/6Ew790f
vqpViqwkS5jKZy40wqyeOAXZttqluKIm6yDrjJ06rLQ35qKZ3UK6agDYlRvkmVe9vUYoTo8sKiB8
kxf95lb10d5hCo2UsKQTD/J8NS9WgwtlUaCEBJqpMjcfv1DXHR7M1iqeF8v9ubjxTTxR0KMsbEms
MaShNUL2y3ujQ/Bfdl5MvSbpS3pnQdzQb7aN4C+I0xhs232qZDAYgnPMGP9ym5hTrNEGT477jJTL
bZEQiOCZsPWMkJAEROCv0bVHtIRlIURgJynBy5N2tfLeVA9pdso/hf1bh+afExb/R+WF94vEOMnY
EGWRBPWOwpQHpZq+/fc2jQX6lpiZ6sP/BIZBNR8Woo3xdtMWBqA3+90Ih/OGxSOdknRRL1wn2Bmv
GIrSJYn6RpY7YF9xm+GaqoGfBD+Lu85kwdLIpBV/Tm0H9pQH2VlrMVEjkp4PcYBsfMBsupDYfN4y
gg4uY45XO6gh7e8i2O2xrbkubIXitVFPGdgaS1w1/GGUC5de/NNkiQOiqma5Mayd34Uq5KpD14nn
y5aDzSkbj26/YnhKOkLKrXI3Zmkwd6Ke6HpdJej2Obqge4oRyCEL3FCqiByru2MLcdyCapL+tYdJ
qC0+IoztQ6TOHYbsTonQObj5dIyzF64m9HURH18sokNPpnmaROjEg7Rr7N238v7IIFWIDwJYDNRM
LnCk8JHkeJrxlv6hYdyrwc4qhOAJbx/NR1wX7pxh5zWCw370xWb7vMUXgWrKIGj9iZlRI6X2b8MU
bgfOkW8c7DscNcec0XqkUKXnlJ5TzMqEesxnEQmmEpzF2gKZivbJ7yxiUE/gfeJiLVyWn4K1VHAS
uo82giF3NUipK0QIlu77B2xakosjqtITLsuC3YtzWKflyC4XSWrYvHxX+rlD/WTesl9WKH3LkS2y
xK/cIVauFZWQTj/2RBiIUPacVX0Bgalahw6SmfWTmWwXsvfJ50OHOWjeVy/3jBEH8bRE4Gg3n3sB
zNPVCpg6Ni9i3TXeeiyt6bTB6u3KmGfOh1zWYwZcQNAwBZjazaN/UZZwMVgbG/yYAI7tO3PNkPBM
r+z97LC+KxpGv25onJU8lWRhyDGbO8Cw4VgHsSae4NZQx6xXsa3DivwUX0Ywf01v8NhHQmPKQZaM
wJe6ly4b8zlnNzXNQ7YBymqGWGAhdcBC/CuPBCIVVIGG1ZhvV4YoUlDx4AsTWtvjE/aObJcIPsZ+
D51jHYHi37CtKoEQaWjv1SdAWsuxtRj7ctvVhNyhjRo/mCw+pY5+XxvIf7s7CHCNSText4ETlGJG
VHjdrweljM+QNFeEWgvfTokCcXx8hMuTZqd7gMa7DokI66Xtf//Jva78bTgXailKAz60rwm2Kw5n
Md3Q+Eua4HGuLO2T2Am08u4vtGlG6B6LExq6Xx8zkxK9QonK+oxPhTzNDxnHhFdZAYUs0tbr5kHA
R+jQxzpBxK8E0KT0YjBtuMNFnkTCAamxckqtm+kf8fcj/47k/tPa28BPle3LQ/fsxEevDB9lZEiD
XBJ0xyzraZbcC51U8vj0cY5p3SFzBSdMYtNd/LsMi1OIFdSNLlXrEHdDLTG92cRLakndTbuPTfOL
lo6DPAgXV6Ro8HEcx3PTYgLzV6m2Hessx9HGYIm5VozShT25meZYWi546z5TB/rJIU4H5woira/U
ittYN3VvNnQBLZgsspW5+tfmiQ59mjTRrkXT4rOU9uxFqGImrcoSLvXd0UmREl5UvKHzvathQ48y
qZS85Eq1I/N9CXL73A7mN7Fe8NJmUWOPZ0RM791N3Zgrq9V6vHlG+qTug7HT+k8PDpbzmDl/8egT
omkIE1zBFQL2gF/0T+LWT+rMXLV5EMmFTmGj1DEO9XdXlFu/LLYAY5B070mmilmg+p1Mmg56/yQt
Q1SzkkZogwOOVZEGStNTifyvaQLV5/yEdTC7S2oblTSy3nE9PUO4kxExgOP7KD8rqh8089Bs0MaQ
/OcqHA5T1zoksOQtd/prBCPCTXlhAGwHWHvkK1+Dh9lLhF2bHtKt1ZzxJYgGVhDIJs6g3TbfGv2+
vACLAu+AfFlF/GXpIK2t7yJd9QFuMseBmfkCfr0F5CLiYb1KbF5amWVPt7LYEKZrJ7Ca7BgegEJM
vfVe3ohf3ktRhtmVLlb+rh7BxYMeEpm0XzWwrTYK2ogUu+QLTeTAaYEDVuXSU/ATlE3qxI8ryWom
X8eREUA6dGEiAqyRkLPGSk9JgKlVleEsJq9TQqKgCd3k6qpFK/MnsVDN09juSO2rWlUNAuIn+gZw
6nk59I4GhZWNEyZtHu+pWsslyqT7fGt89uK8IxZ2l+ax3T0yX9V8Rzkl5hwchAJItqIApB+H81px
SGskQ48LZ8HRgNPADLVoWd3qzNej5OPbQvFXKJ28GcNbGctNPTgEc7ayjjJJ+EYFSaLkvqSFDJxL
TzOs2bq/3tmvgFxkYeyZEYKdepis8f7Qr3s/EU2PR+zPJm2YFKoWb1OM5JVvJno2Xi2ajibzi0AY
IckiEEXHaWducZiRvcIqIQOXtMheD44ZzkrQdGwDRcnI6S3Mkbl0ZNtVNbxyLaN0dZDmgubLlRc0
mJdgQzQt501AP3TyOi+KHD5kOpcDtV9ql5HQh7Ms6Il3yX9octUq0bZolqGmnAXbk2dfIWXwb1r1
961bN2yGXMiWh75oFXnQjDIceFpeOhgJGPd53YPvbPsa5KBQZ45d+VuwTDOzjOW9w0pBFXXI3ZFi
ScvsToJRhxdKBPZ/9N1h3IpD+vTYpogAqbUCFBiD/n05vLw53ApWE7kXBbBjpsZGGLF0IehG+TmI
o+gZdjwWCoXlY+CJBi8lJmGCEViXE2bQd1APacFtdIcvKUtKh0YdxQDH/V4kOwxrdxAr9xeiYVnO
tbQLcoRRzSAMqAulUrWxl3d1QvY7YSTYSnL57t0pNrqEzC+a7jXk0ERXR0VVGIhxyHoygLCFgc8P
tLpD0OyVSNvl1rA+4fUJcbVLHPrlfjEfCI8Po78ZVJc4fJR7Tnlm7TTV12UJ+g6P7ZIoT3vG/Zyk
h6AqldO5sZcDotYByYCi5ZrruZ4ZqMdDGlE7B5CJ8tOkrIiLZTfMYA4r9uGrYOGaK6j1x7+JA71C
xb1a3AOe3+WtEVTNS3q6uq4ukeizpcoh+38lTW2O4RNjEDbMe404jaQLLE87Fh1F7H0U02+ruMAh
+kQ0OOXoNsuC6byw4/hveovcCqHiPLldG4eDV/Ky+bSl/Xwp6nB7ISIl0PCIIZMYF8DmzKMgfDKw
+J0i6QCGZeJ4oHZnfQojdFnBTG7F+odfkgwUQnNHPH9QfBxwj/GnogQFEm9Gj7iIeze+8hYFPTYQ
gEEI6XBoWo8hx/dROcN4u11brF7JkLglayYXcoWp45df+BMaIA+pheMinh6sl2SP91JaPec/OJ7P
OTTfnEoPlx91KHdIF28iNtJUAttXyEw3EGGYxLZxo6DeKmfrsnbAaL4JKXzLciienk4SLzDNyrQv
M7quiJCeQIXep8Ep7IuRxjCeOl2FbVQfQcX1wXHdibCKd5K5fJgGwDq6O+y8/ONsaq0E8h7nvNCF
nIBJz/l+SeBWbEqb98WHBj4pqpKwS0uBK7g2dRCmOjo1sChM1oWCcaV70YPmJQWFhntmpkeOwDlO
1yrqahuvQE10pF/hFiMlzrFpLQcdldgTl3qcyRFlk30FsfJI8SSjRnSquQpeLMcORaFRnymWpjdn
j3/tlQWsAlX8LBsV/1wygL87zEuI1XQ9wJ/FL1hunnqSbMDwd6CAaOGWyMmr1zHJu/NDhBVwZOzj
0d1INY54MzUa+v9DPoWjnup5FfwIWdP5pw8qjr8umf5BmNyxissXeLO9jnXFLAKGjg0p/XMZQxDp
sC/j7alir6pDYyhaJ2g9t7aHTeB3qzcTY7Ew1wWbVGrnEPP8c1nuMHAvTV7717LvYAXhUzKKULt4
q3p8QSBsJwLjNJw3OBTWZAJMlgmRWcYm95V1MrI94DPZtKBMGJxS6rpMpovGEDmTtzF3q7aflaWa
UysZKEgCnzvsntNNG8jumd7Jbc65hRkOPYgoAAU4OxcbaYBVmWieUvOODnJOd3LyVpcfglvW4Bbd
ojaTHpikBr6hFzPa2yItGoDJFefUL8jgf042jRjXmLn2sW6alxmusrFd5SwzNb3b7FozUIww6QYg
bnXCkpRBWVnFSboy62yrRMApXah86lAFpU+Uj0V19iXxobbyq8tLCPB19s/uPQquCPEtmeFeKV+5
CD0zG9b8jU4ymtAvSBPOvulxFEHTq13cZPimMaNigH37uUENgWHGFHK8ypqSA1xjiKQG7vyTQ9fM
wkNeyf+zA2xBCA5Z8xBRZKimsaCs5xrZgS96wF870vK/2XnYEEcZo4xWdjpPdXRmjgvlytmZ9vj9
J94U5c+gTomsOs8O3ivgV4rlY0v9UqbpR3Mx/7ht2AfWHs+sfO5qGz4Dy7F30aCb2UObwR1NEYjx
9MwHenD0AzkZ6n/RBtYyX+rJX8sCVXMPgkWPl2TrzAr9zMUYKkwIgIgZP3MZT34kZn6NB/kkx/L6
npY9bvYX40OiBsvPgVloinFwoY0Mduitg4G4nSq925wne8fggoOtnCKzI7XbSipvaRnNYjKqba8c
Qwhh99sJNS1e2b+YaPN4uIjkNnra9FwS3LXv5+OTt9zyqKyH2xP5sKPcy916mGOHWnl41Tzf0QGT
A8R3ltPwrlBqd6yv5Cgy+/FTC/PimZ3QwM1fq2U/lR5Nzcx4orxOUflSmhYrsXBPqc1uroHyK4J5
NMOSwOo/53tBvK29Brm3ToCeZ9JrgOcyPe4T2xZz2SIBTZcx5sUUedGPU2Y6FcmwtyjXBUtqsTHu
mCTtwa51RKiac1tJGhoV+zt2r678MA5dwQwylBXH3vLqwxsLkS4wG1liVak0n/CqoZtudNHZlU8x
3kY/jGWsqZ2aqgUeiKjilGnOWgM=
`pragma protect end_protected
