entity intruction_decoder is
	port(
		clk : in std_logic
		instruction_word : in std_logic_vector(15 downto 0);
		
		--
		
	);

end entity