module pawc_tb;

pawc_top u_pawc_top(
	.clk    (clk    ),
    .resetn (resetn )
);

endmodule