// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
w0oETvR+QPynX6DYUfEbEHd4tfh0t3Y0tjvI5dIMGKtQvGFpnyPNopknHwyiayTlUn76L1jC4mdf
h7blyMBH7yF47Y1gX41hZuFOX5ExqeKRdwM+qGH22y+nPHmCs6idzIwyNYX0CeAzVvCZexoAf4Ck
FrUQJHqo9muUJhQ3Pp9L4KiW5t/x9n0H8M1op1P/zULlUGiramsTVrbKZVswXnxL5QCvhGyujmi9
9JcbtmqtImEjDhnfh8WM/TqW9L/6gPjP4f5D9XH/zvWcFk9vlO2q1BoVFVlF75AsxoDhpPR0lVrp
LdNAhTVjXaBC07wBCgut01Yz7pZ6E/0kNV+h3Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5760)
2nhl0TiVVw/QIOsqDV4r/4Qptndoms7httzPFrsJD3JHqZdpc7RBqAFOI/skbaJiF7UAWJPYDDdo
sqLkG/PNFV8CrpzGum3M+maFTAkWZ3cm3MdArhkFQrd3jkRSAVIzcpRNq1tozvsnZfgsy0bSffBI
Je2z6Yza5j6Rj8/IKcwuADl8tsaRW38qsBTRnpfDmH+7TGUExCSbDwqSs8vZ9b9C30LHHpeylh6l
AUDG6IH4HHbbDywmuDyskPOqqPrD+046nYZJRwCzI8jbqwQu6l0B9d9unUIKrcvVC+rp+OPJbxz+
NQ/Qt5USzxFG1NmgZ9OHQTZiGkS82BYJKZRLgOJNDx5qxCjxUcdM8460QwILJNticRiwGXNijQ6Z
pwaS2Gh+XbxHI+jqJrSS+PvtE+1Jm9iVfv5YmDvK86x5Ce72aHPAmH06BuIhWQ6YMBRVo2ECGAuh
YeXue+VpoHz/N2A3qzouBDqqJEvyI5bXKGcXSJHVVQsvquXElCav/0qTrHPv+ZsWJEmLquXVmyh+
HmVTCRCN7e7yX4mjYzzy0g7wjLgWHbhbMDip6z65Z+A9/IEE1IUMsPrx2SnSDUzm2LvADy73xcPz
Tprni7o8P6lvgVghDMSyOMwWTqLRAyEGMKz/CQOyfG4llRsO3Zyi5ITj0mNGitZ2ma8zIl6bdN0x
Zt0sPgyPA81pEI/EUY7PuUS1SDEsQ+TtMLpwNZ1FW6E3MTrQc+rl46fFaskrmRlQvo4HlXahlLqb
bPys19QfMp7eMsRSPUk8Vj0g60LVbZGw3qP2Qpo4nFkCXfVRqZ0l0hM9F5rYvd9WRjwQihR0I9ts
aqcRcIWu7L5BbZfdJDcYxRu8zPC0zJCJzzdJfgb/ABS5sPl1AWPtwIvP5WQOmITGNBlwphly85Ou
0AOT6Wj29x2cTjf/KBzvPSGVBkx1GDumbiJmT5bdawAlaLHMj/ZmxskH/iOoMWndgOCGeQkVSGde
m8J3jM6b4oT7u/2ZYSdl5q+IT17hsTE6a8/FRKZPevDeQqZpyH9OU8CcvYs0c7/8odFcXMyrixEL
VV6Odc8O4sxbbuUrJoYQ7ArkvfzQPXAVQS7MnJNHxmXhaNn1ABy3F9DwDSz0kNNMoC6h78x49ev5
FKmf6+zi66hQKM+/BDFRyYpCfhsxnvkVtAjfAztdyPo/77c/3Er4D3XSLK6pPoqmhBavG18+Omhy
nAY0h5dTG+MfrJtou4z5WKc+v+RKQBo++16dafzZGJJ1iMnv6dOkDGnSBPyFYWs6qHAgtjOnrGPh
tWUF96Xn8ZWp/o/Tp/i7md+oI0c3VIiSnN+JxXkd39Xjdg4SW40j9f0SELB0YmTuJ7DbIgE8/ej1
FzhmSpTG4yHgn8HAXEn5QL78mGSGGY1TchqEeG/YkBmTV6AytseNJfA8/3ATbCTBiEuKyZFHViO0
mlyvLu4H6YN9NV6GfJ4ukg9dy3Vf07SLp9VKKVGS5XfU4+EFyvsxJyZA9ahX8gsNEGph1MWAoVte
5x9Ub3FLTBIbtC9feeaG1m8OdoaAungctfUvChw9c2G3TiWTIVBiOMDF6FXORqrk+bv6cBIzlyZ6
SAKESz7U8Qrn6p7/zuKx4oaAXEMiOv1COe+v/NvWLSDN33SlR8b56fQR02bCBUmWGHphlxOmAJ/z
Uurw2PBFb8BlPTggGyX2ywnxX5yk1IG5wFWVZM/KhP4IBhy7lau6N4/1ayqGjUStI/DB+SVJ9UYw
qE/04/nfAeGTyDxkRf3iDs5BmTg+tUPG9Pau1mWrtHNHiOvLg3A3Y6cEEuJ8BIJeA4iQ86ZfyO+i
TFO0tGVA1VWKQ3lbaVRwdUzANqdrg+ePDDB+INaKhRd28rxLkYPzDgxTdHfhfro5Gnrq14F7vyBj
B1RoFvIKOVjyB8uA9LWIfD/T90XHWhgBTS1C0j9OV20kxHbHYgJmBIAMOgPVOW2MNxwuhj6jpra7
DcFMQ4kFihOIl/T+MGI5PZUL0J/DlTUdw+Yi9M2ykFpli2n/+v+Z79Ma6lOHYJXvdFHQ2b7kPM1Y
NTlwQIwcIOW3Jxir3giaxurES1iuZmqFIFs/jRmX0J433HBuOuPPgL3lS4JNRsEtmOy0VcVP7s3Q
NisNIKqqwp1Yge1NOkNE8NY/5S6mvIu7T+e35exSqsMdOK3coez7fMNzCQmyYmZLGPzFkJ81FPOb
AFzJofdLTtSz8kZlBITNiTxpq+YSUCTBeWP3+3xnYqaXiCbUXDBlcIe9ZJwAuUNM9AJHTVDUeAWX
Ihx7panNn3x2UQzcCmTXWr8D7HvbyPaUZLzBldJBELWgPtX3JQSPCv5F/v31upBedYRlXBC3Om1g
mV64CLAb7FXSLtVI6LXSZZ9xwwvRE23BMjJV0T61ICfjgx+s8MuwBy1pYDjfr799jVOMm+rNVoOk
jV8LggL+NsaqBmn1zq8KLpqkRzQdCNbJnWcu/CXl7vLTZO8pbd6MioMUAfsy/gX0IiUbVWbshnF3
w2P1zL73jKzZwjKvLOr9WCofOCVMnrYkdtSFsqfofgb+tiM1LjcdoISkq/9HbRFoGZDWBm9JMASV
4l3zOJQIwWRbY1XJvcwotbQoNxH8cVvnXk+tPKmTXKU8+CxMgD5ZiLIsZXJFWNEBjpzBhRwx5xuo
1KVONkp5u/pk5vu9MpKgc/JOoz0uSlShImfKtMj79Rt/L+3xmYRc0a5dwF+ZcdEond0A1Q2VO344
n5Xj3xPmd/Wb2/EIxKAMXbzq1Fxfbc3P3GdYQf7NvvO56KW8BIdexNfhpGv42eKFTAelTIjAByAp
CDrVyjoCXeNwEL7mFVmHES/CascjagBzrABBFwyEFDQ9AMyVnLi6+WjrvCRkMWidCJGiA8bqzzEz
IMIm5lGv+Zsqnj9fCgKRDRV52aFyYHDq/weL+YJRNRw7qmK801FQ02e64rjwsDxxHEtw2vH61utq
Ee6CfoI2TYPpJriBQoZ8CV7FZ4hj4615cCilgajKblhzTRZmH/ahsaSYQFQak0ctcblC37E+Wa9+
nPmqh1SdGemYh3aVJMbvl+DUNic6OniSF49KKKdP0ayrD42OJ2BA02oC8OUU9UAEIvNg1Ns9Zh9v
5ttOTPDF/ZcjWQ+GMtVjemfGzUnXTYunKKR+2tTjRtdQ3uq+utPebGKMe+TA3099LXGDd0G3J3+0
n72WQjNbqNi3tYN5V0SgPdVqreK0gZgcRYljbYbZipA1BaZ46F6RgF9RNAgkj31AhjqlldtrcCwf
B33eSlOVSs85R9F7Q5XN+6vq3VaAN9fY+nsVAtMk9rueA4qrOvarg7kuBEWXJvj6Ni5zxvhlSao1
HdwpunGV2z2OgXxNBzNHri2m+odJcv7eMHYwuRMEQMQk+t9Dm83cYDupynaNdbKrjdPppRNQiJ1x
obnBj3MKczN1Ci5Fs0YE/2fcsloOqdwAts3PtrnBaOj2nFNszGDg69/ZNLK+wg3//oshTmAhxnjO
g4fx46MPV6qre1oH4HGLWexNaD0R6XfWFT2/VY8Pyoi3Mb/Lbw9w5TIL2/6kIFW2D5vmNQtq3VAp
k+vZJqcOio/8V9x0ZVsb0z1TI5HPnHQ/ys68bVOOpI//FfuTvZAx5egvfgF8qy+S1UNWjDKglARU
DSQbIqd/dP3mYdMp80lk9GKTfmzQ2+RimpUfWytLTOKqR9jgqQoZR1lJrfaGbAqEhaKRh2lmPI9h
/MEmcA4KPm0YM0m+MBKlpnhiQn3HXAHpJIAMFAHKh71vc2XNKomOTtfChinceQf7u9wd5SvBjax3
yr1XhZoevEpNiX0vm45sS++FJFEEXZgkGmaFU2VrGdcuWs/GdtDCagvEaG5zAfmnssT1FtyGomoz
ahppY2LgT+ZFImPQ+gBRP4bIaa8dQ8c2+DD+W//y3IPqPcqZuW0WiwaX3mVY2AopHCNfiBLb6CVL
XpR4PEAOdSj5+tqq7fECLGeFkGTR4n5Hd2a2VUVsZJdrHGGkakb0Bac0pcGm6LHQDIW0e3bG9Xu9
Ltn8sH8KkjAL8T1fSdm+/27VxBRbik06+HB1eui1XoIaEYil9LwSnkE2CnSprcuu3xd7WQ1iLlZP
O91Xv3lSPaxm9X0jdskLajw0m6np4HN7DZPNl1fgyYvR82DLmElbeZ3WnxIqqGTLeYPNEQqNs+sr
JpIvxbTSnEki6QdquaX6+rYb9++ZRnHHIh3Rje+U+1gcDxrXs42xUx9r/UpnA0lUajFDecA1Vbv1
F83Q5rarVzXoQZrUXjoiZpglmgVatM+3lp/RnbReJwboQVMH10C8HBx/pe1tGsGoAVA3olN5QExu
TCidZ/xNexo3sy4ClQFdV4Psm0Y0w1H9b/7wUK9otC8Yfg0Y29dNmmI0kfMsT2LIIIYe9CiMSS4g
5Qx1MKgzUfC1KszQaBw4K27Jfxwe7OyNLX4zFd2ZT+GRILuZKpE/4L+GfHYKhQ/DUpmPoAhH1Pff
hCiqKZxXgPDOAHJ2Fgiak3awYNF8f8+mM/l7RAgOwaM2K/MvWSk3m9AhiPEkF4mg6vNWDAyT9GnE
AT6CpONaEztLxyJkgf7l+FO8NmgmrKJhD1Ul5ejpRsk/AZOLBtWk0mApXJTIYHz1piUfUH25MhEL
Tz7CEC+YxEaFbo8CuqYK1EGBrkHALbpQas/31X2zzSMXZ0kTLy6LS9udBtfwlIUpeX+cz+d9frwK
ggGP5Bvt/no9VWpY9tdlVykyIlG8caFmrNmuH3RhkpVW6793OXf9t8mFC6+NsnB+tbHLcjvSdshE
6SvhsOCpFQrTm+Vd0jWy5Y1MUERFgwlcWFDkng4PxOxzW2ijf261H+kvBFx/OEZLRMzDdoPUsGge
AqBz1+2NXBNeeL40Txl7imW2rDUbC48QWgcZK5S+E73YjwEJW3zQJ1uaTEA3DP/+NHE0sURzWKsk
nFIjucvz3c3MDL7PI4kn1heOvgHuZ0uTpEVIpf4aqj+0OdnNRU2zp60xqHMIiyUfmwepfXo1i+9R
tS1GpjQMqVjpkE+hO6saXArHqV/ArsM2JSCn6FN7NtlzyPyhMxAF3A+mVQxAqdzArPnZoUIRfNl8
uPDsaqMpOkdvdTgnrjJYgAs9hLFuadctnxcC/kTJvbGt7G0ffedoD9SochDfl5QKjBHj1vvorc7v
MSNUxZnJ5OyFHiV+2KmaXUjdOMRUuGlbZC7LVErvBub+nFUPH+O861TK3faAHtt1QNqaNxRrMfzG
oQuVqwXiZDI+DxFMJhg7xXGlKCah5MZzZMKkt5D3nOHTxOY3n5QqYRQesanalwneKcVBLv/tuPO/
fK+SuvUjYwenRLuTllLCsBZJRe5Dbm/L9ZYkhTbJZPeSN7UE+NAeG4ylnKOxhGS317gLvCSZwfYh
cxn1ickYMkjtY6GIQLLYROoj0JbuePRHkuI55x3PCC7up+HZrJT87H3OBHYNA8RPlS0P9Q/PUwQM
3127TMMucr5+9xEBZf1c1lOZxZs4JRSQOa6CIKn1+iadl6CHM+I1Sz1tqao98QtfghlUeqd/MwcK
88Po+3ZE1Dbv+uWEzdkurclvWiIF9C/3qI8Uo7TKhKm/M2hZeEsRBuE9uXklVjjLvZ1ai5UJtiGy
V1yD4RdB+uPVRsHS+adhdktY2vh9XM3hD0lIZSR+3xfVX3ijd5/BdpOZDpOhg4Z5rVQbsvGmynDa
1ZN/2/WpbS9/LMsreAYB3xvGraTm649NqE/CXcQN5nEpnIjz+yEtshYzrA7XSkLiwME2U1a6S9ib
4BF2ZRhyBtr9/0JNDpL4gNjc0sooSB+XqZF8dqTDc9wz3aZFzIHItoDhTqeqkBB6OyZIaG4nQtuE
MNbwddLhsfahh8KE1wLgpYxMRdGxyaV7/uuT1MC4wBbtljT445EI7REQgt6nQR9eVFdrdRf46bI2
OQLC5YE1CzpRAmSXlFuE6m33Zmu08SPBdb4CHSDvoyoSd7VJPWmBDDZuRaFX9Tr3TK8v1UDT80+1
cMUcrwuGONV2g9OEHIkZZ4QYP3xwZ/juSrWX1ODZ/72+M3O93atsEJ1TvMteHPZ+Ww7OeMOwrq7P
ahFWhbZP9vsIYvvRAFxFUxWp7eZpUlz3xLqcXfher7NXUsaKGUjFEl0gIOAowvgRILws5wftGJ//
GW6Gv1Y+perxns6H6JxMGVduqOfVcCAP9ZvT7aE09MtjKVdXYIt4VYx1pCsEAvgIiHBq1U/FRQCT
7SkIpsxDy4PK6AvBQqy9H7aAYaz+8xJo7PMIT2Dlz/QBVS6IdX6Adsmz9nKkCd9gPzErvweyHN2a
vyF1OKaGuQy2oEGR3uX0rRA/J/C7ZMc8IM01KaiZ4W5MKegbc747Q4K0tnZJt3q09qYdNsdFJv1B
HlPZMVcIORHIlvuAOCXRbKL1IgHYl/v+1cA2Reus5wrS/SQjX8DXxTYqs9i/fvUa9KOD0tEbozf9
SMByc0bgNpoO50VI72p9V1q9y4gpqxkHg1AfkFgijlguibMFRbrXMhhbxDLefLY1I60pOxdV6MuI
Jq0DaHYGc1rrIAYcPgPE50WOioQhE7EuqZdBAU46j5L10QinqyzXFTgdlzqlPc+E1UCXvjGGFHeG
2eKAMm3BPabVp19aSppN4gg6ha2SnFhLn3eT92Ytnni2+ua/lNv0T4NZnvYmRV3hq2k1jri6EUdl
OPGrfAbvb4uNa10LO73K6wyP6l+8R1bMBzrptn6g9FwX/1Ol7OSy1Sq/IXy/s68rWjqxlsOsNu91
IfWpSfpmYuC7jJ1HatqQWLi2zBdSPyiMVNa1DaOEP89+hb6/S5+jSbZ2ZVr15AsDjETTduNFT3Gy
BPc/IGqQQQ+M/OFAfQXAGKh7yVfYtuWXJLb4MQlFrT/x6k+ON1zC39VfNwjg+meB+mDYUmZ19lnJ
hyPdMRiKOB1Asiklzgt7VYgQpvmUkP4W4Zx28WS3hR1oTpckPX8ZMDGqO3iTcXgKZqX5FV6+Bxxl
hq6uzPlUgtQdsqm98Kl/T3uieqZs5BofASA4JuZoBKcnjhtGWWgMduoTn+4JK+JGmnGV8GFaseld
Md3BEE5CAlVbvj2hSrt0a/lbo60hwvFDZ18cY6H0DhNNK3LK/1N7WOAWQ9GZQ/kyTZB1XkWaYtnj
CFUgp/TkgdSnzqd+AhscIx16Xzud0+pEfciyBJTKcTfce6NHe4xkACqO5u1DqgZWerkPHGWybNjA
J5t1FQRtLok/ANJm+FvZ+5GtwPM4ESIG3LE3jkVIq0vKqKA+U3HIKYkrCl4i3n/DyTYs/CRlt7CW
qAE0/p13fp95XcmhMbmz3dNedBzSgiTS0lgiFeInrQqjwd9TyFp4brbcgAYraqWjaUvFCw0KFAuu
sI6Id+/6A31sQBWQVds/WDgJEuK4u9ZSU0FZFuLLrwfYWdVHNJ68t7YZiUu5fQ7HMB5cVAsivzvE
5Itc+pHIxrEkVDlY3uLJOHrQqkzA4vkHal/r/gnMMMq78wOKAuNTCP/Bw/5uyVGNJMwHfpB/iAgW
U6a3OK7kNdral62s+thMCg5UD/GevEU/Q/NWd7ELDZH3TBM2X2XqkTN3Nw3QW/drHTX0PimDo51c
P4BlZaMshgx5gFeKax8hhuvLOfLRWKVbzEugWIX8yIjBEgDLOVWpcpmG+GvF6Y97g7f/0UuTGIh5
+4bb
`pragma protect end_protected
