-- WiPhase_top_level_tb.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity WiPhase_top_level_tb is
end entity WiPhase_top_level_tb;

architecture rtl of WiPhase_top_level_tb is
	component WiPhase_top_level is
		port (
			eth_mac_mdio_connection_mdc         : out std_logic;                                       -- mdc
			eth_mac_mdio_connection_mdio_in     : in  std_logic                    := 'X';             -- mdio_in
			eth_mac_mdio_connection_mdio_out    : out std_logic;                                       -- mdio_out
			eth_mac_mdio_connection_mdio_oen    : out std_logic;                                       -- mdio_oen
			eth_mac_rgmii_connection_rgmii_in   : in  std_logic_vector(3 downto 0) := (others => 'X'); -- rgmii_in
			eth_mac_rgmii_connection_rgmii_out  : out std_logic_vector(3 downto 0);                    -- rgmii_out
			eth_mac_rgmii_connection_rx_control : in  std_logic                    := 'X';             -- rx_control
			eth_mac_rgmii_connection_tx_control : out std_logic;                                       -- tx_control
			eth_mac_status_connection_set_10    : in  std_logic                    := 'X';             -- set_10
			eth_mac_status_connection_set_1000  : in  std_logic                    := 'X';             -- set_1000
			eth_mac_status_connection_eth_mode  : out std_logic;                                       -- eth_mode
			eth_mac_status_connection_ena_10    : out std_logic;                                       -- ena_10
			eth_rgmii_rx_clk_clk                : in  std_logic                    := 'X';             -- clk
			eth_rgmii_tx_clk_clk                : in  std_logic                    := 'X';             -- clk
			mclk_i_clk                          : in  std_logic                    := 'X';             -- clk
			mclk_reset_reset_n                  : in  std_logic                    := 'X';             -- reset_n
			pll_inclk_clk                       : in  std_logic                    := 'X';             -- clk
			pll_out_clk                         : out std_logic;                                       -- clk
			sample_pll_areset_conduit_export    : in  std_logic                    := 'X';             -- export
			sample_pll_locked_conduit_export    : out std_logic;                                       -- export
			spi_signals_o_MISO                  : in  std_logic                    := 'X';             -- MISO
			spi_signals_o_MOSI                  : out std_logic;                                       -- MOSI
			spi_signals_o_SCLK                  : out std_logic;                                       -- SCLK
			spi_signals_o_SS_n                  : out std_logic_vector(2 downto 0)                     -- SS_n
		);
	end component WiPhase_top_level;

	component altera_conduit_bfm is
		port (
			sig_mdc      : in  std_logic_vector(0 downto 0) := (others => 'X'); -- mdc
			sig_mdio_in  : out std_logic_vector(0 downto 0);                    -- mdio_in
			sig_mdio_oen : in  std_logic_vector(0 downto 0) := (others => 'X'); -- mdio_oen
			sig_mdio_out : in  std_logic_vector(0 downto 0) := (others => 'X')  -- mdio_out
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			sig_rgmii_in   : out std_logic_vector(3 downto 0);                    -- rgmii_in
			sig_rgmii_out  : in  std_logic_vector(3 downto 0) := (others => 'X'); -- rgmii_out
			sig_rx_control : out std_logic_vector(0 downto 0);                    -- rx_control
			sig_tx_control : in  std_logic_vector(0 downto 0) := (others => 'X')  -- tx_control
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			sig_ena_10   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- ena_10
			sig_eth_mode : in  std_logic_vector(0 downto 0) := (others => 'X'); -- eth_mode
			sig_set_10   : out std_logic_vector(0 downto 0);                    -- set_10
			sig_set_1000 : out std_logic_vector(0 downto 0)                     -- set_1000
		);
	end component altera_conduit_bfm_0003;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm_0004 is
		port (
			sig_export : out std_logic_vector(0 downto 0)   -- export
		);
	end component altera_conduit_bfm_0004;

	component altera_conduit_bfm_0005 is
		port (
			sig_export : in std_logic_vector(0 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0005;

	component altera_conduit_bfm_0006 is
		port (
			sig_MISO : out std_logic_vector(0 downto 0);                    -- MISO
			sig_MOSI : in  std_logic_vector(0 downto 0) := (others => 'X'); -- MOSI
			sig_SCLK : in  std_logic_vector(0 downto 0) := (others => 'X'); -- SCLK
			sig_SS_n : in  std_logic_vector(2 downto 0) := (others => 'X')  -- SS_n
		);
	end component altera_conduit_bfm_0006;

	signal wiphase_top_level_inst_eth_rgmii_rx_clk_bfm_clk_clk                    : std_logic;                    -- WiPhase_top_level_inst_eth_rgmii_rx_clk_bfm:clk -> [WiPhase_top_level_inst:eth_rgmii_rx_clk_clk, WiPhase_top_level_inst_mclk_reset_bfm:clk]
	signal wiphase_top_level_inst_eth_rgmii_tx_clk_bfm_clk_clk                    : std_logic;                    -- WiPhase_top_level_inst_eth_rgmii_tx_clk_bfm:clk -> WiPhase_top_level_inst:eth_rgmii_tx_clk_clk
	signal wiphase_top_level_inst_mclk_i_bfm_clk_clk                              : std_logic;                    -- WiPhase_top_level_inst_mclk_i_bfm:clk -> WiPhase_top_level_inst:mclk_i_clk
	signal wiphase_top_level_inst_pll_inclk_bfm_clk_clk                           : std_logic;                    -- WiPhase_top_level_inst_pll_inclk_bfm:clk -> WiPhase_top_level_inst:pll_inclk_clk
	signal wiphase_top_level_inst_eth_mac_mdio_connection_bfm_conduit_mdio_in     : std_logic_vector(0 downto 0); -- WiPhase_top_level_inst_eth_mac_mdio_connection_bfm:sig_mdio_in -> WiPhase_top_level_inst:eth_mac_mdio_connection_mdio_in
	signal wiphase_top_level_inst_eth_mac_mdio_connection_mdio_oen                : std_logic;                    -- WiPhase_top_level_inst:eth_mac_mdio_connection_mdio_oen -> WiPhase_top_level_inst_eth_mac_mdio_connection_bfm:sig_mdio_oen
	signal wiphase_top_level_inst_eth_mac_mdio_connection_mdio_out                : std_logic;                    -- WiPhase_top_level_inst:eth_mac_mdio_connection_mdio_out -> WiPhase_top_level_inst_eth_mac_mdio_connection_bfm:sig_mdio_out
	signal wiphase_top_level_inst_eth_mac_mdio_connection_mdc                     : std_logic;                    -- WiPhase_top_level_inst:eth_mac_mdio_connection_mdc -> WiPhase_top_level_inst_eth_mac_mdio_connection_bfm:sig_mdc
	signal wiphase_top_level_inst_eth_mac_rgmii_connection_tx_control             : std_logic;                    -- WiPhase_top_level_inst:eth_mac_rgmii_connection_tx_control -> WiPhase_top_level_inst_eth_mac_rgmii_connection_bfm:sig_tx_control
	signal wiphase_top_level_inst_eth_mac_rgmii_connection_bfm_conduit_rx_control : std_logic_vector(0 downto 0); -- WiPhase_top_level_inst_eth_mac_rgmii_connection_bfm:sig_rx_control -> WiPhase_top_level_inst:eth_mac_rgmii_connection_rx_control
	signal wiphase_top_level_inst_eth_mac_rgmii_connection_bfm_conduit_rgmii_in   : std_logic_vector(3 downto 0); -- WiPhase_top_level_inst_eth_mac_rgmii_connection_bfm:sig_rgmii_in -> WiPhase_top_level_inst:eth_mac_rgmii_connection_rgmii_in
	signal wiphase_top_level_inst_eth_mac_rgmii_connection_rgmii_out              : std_logic_vector(3 downto 0); -- WiPhase_top_level_inst:eth_mac_rgmii_connection_rgmii_out -> WiPhase_top_level_inst_eth_mac_rgmii_connection_bfm:sig_rgmii_out
	signal wiphase_top_level_inst_eth_mac_status_connection_ena_10                : std_logic;                    -- WiPhase_top_level_inst:eth_mac_status_connection_ena_10 -> WiPhase_top_level_inst_eth_mac_status_connection_bfm:sig_ena_10
	signal wiphase_top_level_inst_eth_mac_status_connection_eth_mode              : std_logic;                    -- WiPhase_top_level_inst:eth_mac_status_connection_eth_mode -> WiPhase_top_level_inst_eth_mac_status_connection_bfm:sig_eth_mode
	signal wiphase_top_level_inst_eth_mac_status_connection_bfm_conduit_set_1000  : std_logic_vector(0 downto 0); -- WiPhase_top_level_inst_eth_mac_status_connection_bfm:sig_set_1000 -> WiPhase_top_level_inst:eth_mac_status_connection_set_1000
	signal wiphase_top_level_inst_eth_mac_status_connection_bfm_conduit_set_10    : std_logic_vector(0 downto 0); -- WiPhase_top_level_inst_eth_mac_status_connection_bfm:sig_set_10 -> WiPhase_top_level_inst:eth_mac_status_connection_set_10
	signal wiphase_top_level_inst_sample_pll_areset_conduit_bfm_conduit_export    : std_logic_vector(0 downto 0); -- WiPhase_top_level_inst_sample_pll_areset_conduit_bfm:sig_export -> WiPhase_top_level_inst:sample_pll_areset_conduit_export
	signal wiphase_top_level_inst_sample_pll_locked_conduit_export                : std_logic;                    -- WiPhase_top_level_inst:sample_pll_locked_conduit_export -> WiPhase_top_level_inst_sample_pll_locked_conduit_bfm:sig_export
	signal wiphase_top_level_inst_spi_signals_o_sclk                              : std_logic;                    -- WiPhase_top_level_inst:spi_signals_o_SCLK -> WiPhase_top_level_inst_spi_signals_o_bfm:sig_SCLK
	signal wiphase_top_level_inst_spi_signals_o_ss_n                              : std_logic_vector(2 downto 0); -- WiPhase_top_level_inst:spi_signals_o_SS_n -> WiPhase_top_level_inst_spi_signals_o_bfm:sig_SS_n
	signal wiphase_top_level_inst_spi_signals_o_bfm_conduit_miso                  : std_logic_vector(0 downto 0); -- WiPhase_top_level_inst_spi_signals_o_bfm:sig_MISO -> WiPhase_top_level_inst:spi_signals_o_MISO
	signal wiphase_top_level_inst_spi_signals_o_mosi                              : std_logic;                    -- WiPhase_top_level_inst:spi_signals_o_MOSI -> WiPhase_top_level_inst_spi_signals_o_bfm:sig_MOSI
	signal wiphase_top_level_inst_mclk_reset_bfm_reset_reset                      : std_logic;                    -- WiPhase_top_level_inst_mclk_reset_bfm:reset -> WiPhase_top_level_inst:mclk_reset_reset_n

begin

	wiphase_top_level_inst : component WiPhase_top_level
		port map (
			eth_mac_mdio_connection_mdc         => wiphase_top_level_inst_eth_mac_mdio_connection_mdc,                        --   eth_mac_mdio_connection.mdc
			eth_mac_mdio_connection_mdio_in     => wiphase_top_level_inst_eth_mac_mdio_connection_bfm_conduit_mdio_in(0),     --                          .mdio_in
			eth_mac_mdio_connection_mdio_out    => wiphase_top_level_inst_eth_mac_mdio_connection_mdio_out,                   --                          .mdio_out
			eth_mac_mdio_connection_mdio_oen    => wiphase_top_level_inst_eth_mac_mdio_connection_mdio_oen,                   --                          .mdio_oen
			eth_mac_rgmii_connection_rgmii_in   => wiphase_top_level_inst_eth_mac_rgmii_connection_bfm_conduit_rgmii_in,      --  eth_mac_rgmii_connection.rgmii_in
			eth_mac_rgmii_connection_rgmii_out  => wiphase_top_level_inst_eth_mac_rgmii_connection_rgmii_out,                 --                          .rgmii_out
			eth_mac_rgmii_connection_rx_control => wiphase_top_level_inst_eth_mac_rgmii_connection_bfm_conduit_rx_control(0), --                          .rx_control
			eth_mac_rgmii_connection_tx_control => wiphase_top_level_inst_eth_mac_rgmii_connection_tx_control,                --                          .tx_control
			eth_mac_status_connection_set_10    => wiphase_top_level_inst_eth_mac_status_connection_bfm_conduit_set_10(0),    -- eth_mac_status_connection.set_10
			eth_mac_status_connection_set_1000  => wiphase_top_level_inst_eth_mac_status_connection_bfm_conduit_set_1000(0),  --                          .set_1000
			eth_mac_status_connection_eth_mode  => wiphase_top_level_inst_eth_mac_status_connection_eth_mode,                 --                          .eth_mode
			eth_mac_status_connection_ena_10    => wiphase_top_level_inst_eth_mac_status_connection_ena_10,                   --                          .ena_10
			eth_rgmii_rx_clk_clk                => wiphase_top_level_inst_eth_rgmii_rx_clk_bfm_clk_clk,                       --          eth_rgmii_rx_clk.clk
			eth_rgmii_tx_clk_clk                => wiphase_top_level_inst_eth_rgmii_tx_clk_bfm_clk_clk,                       --          eth_rgmii_tx_clk.clk
			mclk_i_clk                          => wiphase_top_level_inst_mclk_i_bfm_clk_clk,                                 --                    mclk_i.clk
			mclk_reset_reset_n                  => wiphase_top_level_inst_mclk_reset_bfm_reset_reset,                         --                mclk_reset.reset_n
			pll_inclk_clk                       => wiphase_top_level_inst_pll_inclk_bfm_clk_clk,                              --                 pll_inclk.clk
			pll_out_clk                         => open,                                                                      --                   pll_out.clk
			sample_pll_areset_conduit_export    => wiphase_top_level_inst_sample_pll_areset_conduit_bfm_conduit_export(0),    -- sample_pll_areset_conduit.export
			sample_pll_locked_conduit_export    => wiphase_top_level_inst_sample_pll_locked_conduit_export,                   -- sample_pll_locked_conduit.export
			spi_signals_o_MISO                  => wiphase_top_level_inst_spi_signals_o_bfm_conduit_miso(0),                  --             spi_signals_o.MISO
			spi_signals_o_MOSI                  => wiphase_top_level_inst_spi_signals_o_mosi,                                 --                          .MOSI
			spi_signals_o_SCLK                  => wiphase_top_level_inst_spi_signals_o_sclk,                                 --                          .SCLK
			spi_signals_o_SS_n                  => wiphase_top_level_inst_spi_signals_o_ss_n                                  --                          .SS_n
		);

	wiphase_top_level_inst_eth_mac_mdio_connection_bfm : component altera_conduit_bfm
		port map (
			sig_mdc(0)      => wiphase_top_level_inst_eth_mac_mdio_connection_mdc,                 -- conduit.mdc
			sig_mdio_in     => wiphase_top_level_inst_eth_mac_mdio_connection_bfm_conduit_mdio_in, --        .mdio_in
			sig_mdio_oen(0) => wiphase_top_level_inst_eth_mac_mdio_connection_mdio_oen,            --        .mdio_oen
			sig_mdio_out(0) => wiphase_top_level_inst_eth_mac_mdio_connection_mdio_out             --        .mdio_out
		);

	wiphase_top_level_inst_eth_mac_rgmii_connection_bfm : component altera_conduit_bfm_0002
		port map (
			sig_rgmii_in      => wiphase_top_level_inst_eth_mac_rgmii_connection_bfm_conduit_rgmii_in,   -- conduit.rgmii_in
			sig_rgmii_out     => wiphase_top_level_inst_eth_mac_rgmii_connection_rgmii_out,              --        .rgmii_out
			sig_rx_control    => wiphase_top_level_inst_eth_mac_rgmii_connection_bfm_conduit_rx_control, --        .rx_control
			sig_tx_control(0) => wiphase_top_level_inst_eth_mac_rgmii_connection_tx_control              --        .tx_control
		);

	wiphase_top_level_inst_eth_mac_status_connection_bfm : component altera_conduit_bfm_0003
		port map (
			sig_ena_10(0)   => wiphase_top_level_inst_eth_mac_status_connection_ena_10,               -- conduit.ena_10
			sig_eth_mode(0) => wiphase_top_level_inst_eth_mac_status_connection_eth_mode,             --        .eth_mode
			sig_set_10      => wiphase_top_level_inst_eth_mac_status_connection_bfm_conduit_set_10,   --        .set_10
			sig_set_1000    => wiphase_top_level_inst_eth_mac_status_connection_bfm_conduit_set_1000  --        .set_1000
		);

	wiphase_top_level_inst_eth_rgmii_rx_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => wiphase_top_level_inst_eth_rgmii_rx_clk_bfm_clk_clk  -- clk.clk
		);

	wiphase_top_level_inst_eth_rgmii_tx_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => wiphase_top_level_inst_eth_rgmii_tx_clk_bfm_clk_clk  -- clk.clk
		);

	wiphase_top_level_inst_mclk_i_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => wiphase_top_level_inst_mclk_i_bfm_clk_clk  -- clk.clk
		);

	wiphase_top_level_inst_mclk_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => wiphase_top_level_inst_mclk_reset_bfm_reset_reset,   -- reset.reset_n
			clk   => wiphase_top_level_inst_eth_rgmii_rx_clk_bfm_clk_clk  --   clk.clk
		);

	wiphase_top_level_inst_pll_inclk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => wiphase_top_level_inst_pll_inclk_bfm_clk_clk  -- clk.clk
		);

	wiphase_top_level_inst_sample_pll_areset_conduit_bfm : component altera_conduit_bfm_0004
		port map (
			sig_export => wiphase_top_level_inst_sample_pll_areset_conduit_bfm_conduit_export  -- conduit.export
		);

	wiphase_top_level_inst_sample_pll_locked_conduit_bfm : component altera_conduit_bfm_0005
		port map (
			sig_export(0) => wiphase_top_level_inst_sample_pll_locked_conduit_export  -- conduit.export
		);

	wiphase_top_level_inst_spi_signals_o_bfm : component altera_conduit_bfm_0006
		port map (
			sig_MISO    => wiphase_top_level_inst_spi_signals_o_bfm_conduit_miso, -- conduit.MISO
			sig_MOSI(0) => wiphase_top_level_inst_spi_signals_o_mosi,             --        .MOSI
			sig_SCLK(0) => wiphase_top_level_inst_spi_signals_o_sclk,             --        .SCLK
			sig_SS_n    => wiphase_top_level_inst_spi_signals_o_ss_n              --        .SS_n
		);

end architecture rtl; -- of WiPhase_top_level_tb
